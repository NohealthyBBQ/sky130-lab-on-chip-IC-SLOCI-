magic
tech sky130A
timestamp 1662864467
<< locali >>
rect -8750 6930 17690 6960
<< metal1 >>
rect -8750 7400 17700 7450
rect -8750 6510 -8700 7400
rect 17650 6510 17700 7400
rect -8750 6470 17700 6510
rect -8750 4750 -8700 6470
rect 17650 4750 17700 6470
rect -8750 4710 17700 4750
rect -8750 -890 -8700 4710
rect 150 2710 210 2870
rect 1030 2820 1090 2870
rect 1030 2760 1300 2820
rect 2140 2760 2400 2820
rect 3240 2760 3500 2820
rect 4340 2760 4600 2820
rect 5440 2760 5700 2820
rect 6540 2760 6800 2820
rect 7640 2760 7900 2820
rect 1030 2710 1090 2760
rect 370 960 420 1100
rect 830 970 880 1110
rect 1040 1010 1310 1060
rect 2130 1010 2400 1060
rect 3230 1010 3500 1060
rect 4340 1010 4610 1060
rect 5440 1010 5710 1060
rect 6530 1010 6800 1060
rect 7640 1010 7910 1060
rect 17650 -890 17700 4710
rect -8750 -930 17700 -890
rect -8750 -2650 -8700 -930
rect 17650 -2650 17700 -930
rect -8750 -2690 17700 -2650
rect -8750 -3600 -8700 -2690
rect 17650 -3600 17700 -2690
rect -8750 -3650 17700 -3600
use XM_output_mirr_combined  XM_output_mirr_combined_0
timestamp 1662815693
transform 1 0 0 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_1
timestamp 1662815693
transform 1 0 0 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_2
timestamp 1662815693
transform 1 0 0 0 1 -3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_3
timestamp 1662815693
transform 1 0 -8800 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_4
timestamp 1662815693
transform 1 0 -8800 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_5
timestamp 1662815693
transform 1 0 -8800 0 1 -3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_6
timestamp 1662815693
transform 1 0 8800 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_7
timestamp 1662815693
transform 1 0 8800 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_8
timestamp 1662815693
transform 1 0 8800 0 1 -3700
box 0 0 8950 3800
<< labels >>
flabel space 40 44 8913 3752 0 FreeSans 6400 0 0 0 inner_core
<< end >>
