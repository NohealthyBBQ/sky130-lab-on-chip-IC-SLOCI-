magic
tech sky130A
magscale 1 2
timestamp 1661820354
<< metal1 >>
rect 539 2933 549 3013
rect 629 2933 639 3013
rect 1455 2933 1465 3013
rect 1545 2933 1555 3013
rect 2371 2933 2381 3013
rect 2461 2933 2471 3013
rect 81 2425 91 2505
rect 171 2425 181 2505
rect 997 2425 1007 2505
rect 1087 2425 1097 2505
rect 1913 2425 1923 2505
rect 2003 2425 2013 2505
rect 527 2347 617 2393
rect 985 2347 1075 2393
rect 1443 2347 1533 2393
rect 1901 2347 1991 2393
rect 527 1591 617 1637
rect 985 1591 1075 1637
rect 1443 1591 1533 1637
rect 1901 1591 1991 1637
rect 527 835 617 881
rect 985 835 1075 881
rect 1443 835 1533 881
rect 1901 835 1991 881
rect 527 79 617 125
rect 985 79 1075 125
rect 1443 79 1533 125
rect 1901 79 1991 125
<< via1 >>
rect 549 2933 629 3013
rect 1465 2933 1545 3013
rect 2381 2933 2461 3013
rect 91 2425 171 2505
rect 1007 2425 1087 2505
rect 1923 2425 2003 2505
<< metal2 >>
rect 549 3013 629 3023
rect 549 2923 629 2933
rect 1465 3013 1545 3023
rect 1465 2923 1545 2933
rect 2381 3013 2461 3023
rect 2381 2923 2461 2933
rect 91 2505 171 2515
rect 91 2415 171 2425
rect 1007 2505 1087 2515
rect 1007 2415 1087 2425
rect 1923 2505 2003 2515
rect 1923 2415 2003 2425
use sky130_fd_pr__nfet_01v8_USQY94  sky130_fd_pr__nfet_01v8_USQY94_0
timestamp 1661796674
transform 1 0 1259 0 1 1560
box -1312 -1613 1312 1613
<< end >>
