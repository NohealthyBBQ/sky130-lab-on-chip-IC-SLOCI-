magic
tech sky130A
magscale 1 2
timestamp 1662832237
<< nwell >>
rect -8726 10225 -8100 11452
<< locali >>
rect -9000 8140 -8880 8440
<< metal1 >>
rect -10090 8240 -10080 8300
rect -10020 8240 -10010 8300
rect -10080 7780 -9980 7920
<< via1 >>
rect -10080 8240 -10020 8300
<< metal2 >>
rect -10080 8300 -10020 9160
rect -10080 8230 -10020 8240
rect -14220 2430 -14130 2464
use XM_Rref  XM_Rref_0
timestamp 1662826901
transform 0 1 -13057 -1 0 -5305
box -1417 -1173 5029 21223
use XM_bjt  XM_bjt_0
timestamp 1662737136
transform 1 0 -1980 0 1 -2620
box 0 0 6492 9068
use XM_bjt_out  XM_bjt_out_0
timestamp 1662830870
transform 1 0 -1980 0 1 6780
box 0 0 6492 3916
use XM_feedbackmir2  XM_feedbackmir2_0
timestamp 1662719914
transform 1 0 -10781 0 1 9846
box -140 -160 2080 1600
use XM_feedbackmir  XM_feedbackmir_0
timestamp 1662675866
transform 1 0 -13500 0 1 8386
box -700 -500 2900 3100
use XM_otabias_nmos  XM_otabias_nmos_0
timestamp 1662818991
transform 1 0 -10166 0 1 7710
box -53 -53 1339 1105
use XM_otabias_pmos  XM_otabias_pmos_0
timestamp 1662818872
transform 1 0 -10817 0 1 8939
box -53 -53 1571 879
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662816987
transform 1 0 26563 0 1 -3003
box -17600 -7400 35500 15000
use XM_pdn  XM_pdn_0
timestamp 1662820526
transform 1 0 -8791 0 1 9133
box -53 -718 5502 1206
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662739988
transform 1 0 -8840 0 1 1874
box -5380 594 6776 6403
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_1
timestamp 1662739988
transform 1 0 -8840 0 1 -4044
box -5380 594 6776 6403
use sky130_fd_pr__res_high_po_1p41_6ZUZ5C  sky130_fd_pr__res_high_po_1p41_6ZUZ5C_0
timestamp 1662820359
transform 1 0 -8623 0 1 7103
box -307 -1408 307 1408
use sky130_fd_pr__res_high_po_1p41_GWJZ59  sky130_fd_pr__res_high_po_1p41_GWJZ59_0
timestamp 1662827202
transform 0 1 -3232 -1 0 -3669
box -307 -10998 307 10998
use sky130_fd_pr__res_high_po_1p41_HX7ZEK  sky130_fd_pr__res_high_po_1p41_HX7ZEK_0
timestamp 1662827686
transform 0 1 3187 -1 0 -3015
box -307 -5348 307 5348
use sky130_fd_pr__res_high_po_1p41_S8KB58  sky130_fd_pr__res_high_po_1p41_S8KB58_0
timestamp 1662758895
transform 0 1 -3253 -1 0 11177
box -307 -4837 307 4837
<< end >>
