magic
tech sky130A
magscale 1 2
timestamp 1662486559
<< error_s >>
rect 56763 20989 56798 21023
rect 56764 20970 56798 20989
rect 822 15750 1566 15752
rect 822 14954 1566 14956
rect 7798 14799 7833 14833
rect 7799 14780 7833 14799
rect 822 14158 1566 14160
rect 822 13362 1566 13364
rect 3738 12781 3773 12815
rect 3739 12762 3773 12781
rect 822 12566 1566 12568
rect 822 11770 1566 11772
rect 822 10974 1566 10976
rect 822 10178 1566 10180
rect 822 9382 1566 9384
rect 822 8586 1566 8588
rect 822 7790 1566 7792
rect 822 6994 1566 6996
rect 822 6198 1566 6200
rect 822 5402 1566 5404
rect 822 4606 1566 4608
rect 822 3810 1566 3812
rect 822 3014 1566 3016
rect 822 2218 1566 2220
rect 1521 1931 1566 1985
rect 2714 1967 2748 1985
rect 1541 1424 1566 1931
rect 822 1422 1566 1424
rect 1575 1897 1620 1931
rect 822 626 824 1370
rect 1541 626 1566 1370
rect 1575 626 1609 1897
rect 1575 592 1600 626
rect 2678 583 2748 1967
rect 2678 547 2731 583
rect 3219 530 3234 5020
rect 3253 530 3287 5074
rect 3253 496 3268 530
rect 3758 477 3773 12762
rect 3792 12728 3827 12762
rect 4277 12728 4312 12762
rect 3792 477 3826 12728
rect 4278 12709 4312 12728
rect 3792 443 3807 477
rect 4297 424 4312 12709
rect 4331 12675 4366 12709
rect 4331 424 4365 12675
rect 6520 2541 6555 2575
rect 7113 2558 7147 2576
rect 6521 2522 6555 2541
rect 4786 978 4887 1232
rect 5040 488 5141 978
rect 5623 901 5657 920
rect 6035 902 6069 920
rect 5612 866 5657 901
rect 4331 390 4346 424
rect 5632 361 5657 866
rect 5666 832 5711 866
rect 5666 361 5700 832
rect 5812 764 5870 770
rect 5812 730 5824 764
rect 5812 724 5870 730
rect 5812 454 5870 460
rect 5812 420 5824 454
rect 5812 414 5870 420
rect 5666 327 5691 361
rect 5999 318 6069 902
rect 5999 282 6052 318
rect 6540 265 6555 2522
rect 6574 2488 6609 2522
rect 6574 265 6608 2488
rect 6574 231 6589 265
rect 7077 212 7147 2558
rect 7077 176 7130 212
rect 7818 159 7833 14780
rect 7852 14746 7887 14780
rect 7852 159 7886 14746
rect 10752 14481 10787 14515
rect 10753 14462 10787 14481
rect 10067 696 10101 714
rect 9106 664 9164 670
rect 8538 601 8572 655
rect 8960 637 8994 655
rect 7852 125 7867 159
rect 8557 106 8572 601
rect 8591 567 8626 601
rect 8591 106 8625 567
rect 8737 499 8795 505
rect 8737 465 8749 499
rect 8737 459 8795 465
rect 8737 189 8795 195
rect 8737 155 8749 189
rect 8737 149 8795 155
rect 8591 72 8606 106
rect 8924 53 8994 637
rect 9106 630 9118 664
rect 9106 624 9164 630
rect 9844 558 9902 564
rect 9276 531 9310 549
rect 9698 531 9732 549
rect 9276 495 9346 531
rect 9293 461 9364 495
rect 9106 136 9164 142
rect 9106 102 9118 136
rect 9106 96 9164 102
rect 8924 17 8977 53
rect 9293 0 9363 461
rect 9475 393 9533 399
rect 9475 359 9487 393
rect 9475 353 9533 359
rect 9475 83 9533 89
rect 9475 49 9487 83
rect 9475 43 9533 49
rect 9293 -36 9346 0
rect 9662 -53 9732 531
rect 9844 524 9856 558
rect 9844 518 9902 524
rect 9844 30 9902 36
rect 9844 -4 9856 30
rect 9844 -10 9902 -4
rect 9662 -89 9715 -53
rect 10031 -106 10101 696
rect 10031 -142 10084 -106
rect 10772 -159 10787 14462
rect 10806 14428 10841 14462
rect 11491 14428 11526 14462
rect 10806 -159 10840 14428
rect 11492 14409 11526 14428
rect 10806 -193 10821 -159
rect 11511 -212 11526 14409
rect 11545 14375 11580 14409
rect 12230 14375 12265 14409
rect 11545 -212 11579 14375
rect 12231 14356 12265 14375
rect 11545 -246 11560 -212
rect 12250 -265 12265 14356
rect 12284 14322 12319 14356
rect 12284 -265 12318 14322
rect 17207 14269 17242 14303
rect 17208 14250 17242 14269
rect 12284 -299 12299 -265
rect 17227 -371 17242 14250
rect 17261 14216 17296 14250
rect 17261 -371 17295 14216
rect 50165 14163 50200 14197
rect 50166 14144 50200 14163
rect 17261 -405 17276 -371
rect 50185 -477 50200 14144
rect 50219 14110 50254 14144
rect 50904 14110 50939 14144
rect 50219 -477 50253 14110
rect 50905 14091 50939 14110
rect 50219 -511 50234 -477
rect 50924 -530 50939 14091
rect 50958 14057 50993 14091
rect 51643 14057 51678 14091
rect 50958 -530 50992 14057
rect 51644 14038 51678 14057
rect 50958 -564 50973 -530
rect 51663 -583 51678 14038
rect 51697 14004 51732 14038
rect 52382 14004 52417 14038
rect 51697 -583 51731 14004
rect 52383 13985 52417 14004
rect 51697 -617 51712 -583
rect 52402 -636 52417 13985
rect 52436 13951 52471 13985
rect 53121 13951 53156 13985
rect 52436 -636 52470 13951
rect 53122 13932 53156 13951
rect 52436 -670 52451 -636
rect 53141 -689 53156 13932
rect 53175 13898 53210 13932
rect 53860 13898 53895 13932
rect 53175 -689 53209 13898
rect 53861 13879 53895 13898
rect 53175 -723 53190 -689
rect 53880 -742 53895 13879
rect 53914 13845 53949 13879
rect 54599 13845 54634 13879
rect 53914 -742 53948 13845
rect 54600 13826 54634 13845
rect 53914 -776 53929 -742
rect 54619 -795 54634 13826
rect 54653 13792 54688 13826
rect 54653 -795 54687 13792
rect 54653 -829 54668 -795
rect 55358 -848 55373 13826
rect 55392 -848 55426 13880
rect 55392 -882 55407 -848
rect 56783 -901 56798 20970
rect 56817 20936 56852 20970
rect 58188 20936 58223 20970
rect 56817 -901 56851 20936
rect 58189 20917 58223 20936
rect 56817 -935 56832 -901
rect 58208 -954 58223 20917
rect 58242 20883 58277 20917
rect 59613 20883 59648 20917
rect 58242 -954 58276 20883
rect 59614 20864 59648 20883
rect 58242 -988 58257 -954
rect 59633 -1007 59648 20864
rect 59667 20830 59702 20864
rect 61038 20830 61073 20864
rect 59667 -1007 59701 20830
rect 61039 20811 61073 20830
rect 59667 -1041 59682 -1007
rect 61058 -1060 61073 20811
rect 61092 20777 61127 20811
rect 61092 -1060 61126 20777
rect 61092 -1094 61107 -1060
rect 62483 -1113 62498 20811
rect 62517 -1113 62551 20865
rect 63025 8383 63059 8437
rect 62517 -1147 62532 -1113
rect 63044 -1166 63059 8383
rect 63078 8349 63113 8383
rect 63078 -1166 63112 8349
rect 63586 1472 63620 1526
rect 63078 -1200 63093 -1166
rect 63605 -1219 63620 1472
rect 63639 1438 63674 1472
rect 63639 -1219 63673 1438
rect 63639 -1253 63654 -1219
rect 64166 -1272 64181 1472
rect 64200 -1272 64234 1526
rect 64200 -1306 64215 -1272
use sky130_fd_pr__cap_mim_m3_1_ZQCY8R  XC_porst
timestamp 1662486269
transform 1 0 14790 0 1 1746
box -1750 -2100 1749 2100
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM4
timestamp 1662486269
transform 1 0 7473 0 1 7496
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM5
timestamp 1662486269
transform 1 0 8212 0 1 7443
box -396 -7373 396 7373
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM8
timestamp 1662486269
transform 1 0 6834 0 1 1367
box -296 -1191 296 1191
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM11
timestamp 1662486269
transform 1 0 6295 0 1 1420
box -296 -1191 296 1191
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM15
timestamp 1662486269
transform 1 0 10427 0 1 7178
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM16
timestamp 1662486269
transform 1 0 11166 0 1 7125
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM17
timestamp 1662486269
transform 1 0 11905 0 1 7072
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM18
timestamp 1662486269
transform 1 0 12644 0 1 7019
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM19
timestamp 1662486269
transform 1 0 16882 0 1 6966
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM20
timestamp 1662486269
transform 1 0 17621 0 1 6913
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM21
timestamp 1662486269
transform 1 0 49840 0 1 6860
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM22
timestamp 1662486269
transform 1 0 50579 0 1 6807
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM23
timestamp 1662486269
transform 1 0 51318 0 1 6754
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM24
timestamp 1662486269
transform 1 0 52057 0 1 6701
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM25
timestamp 1662486269
transform 1 0 52796 0 1 6648
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM26
timestamp 1662486269
transform 1 0 53535 0 1 6595
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM27
timestamp 1662486269
transform 1 0 54274 0 1 6542
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM28
timestamp 1662486269
transform 1 0 55013 0 1 6489
box -396 -7373 396 7373
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir1
timestamp 1662486269
transform 1 0 4052 0 1 6593
box -296 -6205 296 6205
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir2
timestamp 1662486269
transform 1 0 4591 0 1 6540
box -296 -6205 296 6205
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir
timestamp 1662486269
transform 1 0 3513 0 1 6646
box -296 -6205 296 6205
use sky130_fd_pr__nfet_01v8_648S5X  XMinv_n1
timestamp 1662486269
transform 1 0 9504 0 1 221
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XMinv_n
timestamp 1662486269
transform 1 0 8766 0 1 327
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XMinv_p1
timestamp 1662486269
transform 1 0 9873 0 1 277
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XMinv_p
timestamp 1662486269
transform 1 0 9135 0 1 383
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_lvt_AHZKRZ  XMota_bias_n
timestamp 1662486269
transform 1 0 2135 0 1 1257
box -596 -710 596 710
use sky130_fd_pr__pfet_01v8_lvt_AH4MH9  XMota_bias_p
timestamp 1662486269
transform 1 0 2974 0 1 2775
box -296 -2281 296 2281
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XMpdn
timestamp 1662486269
transform 1 0 5841 0 1 592
box -211 -310 211 310
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 0 796 0 33 796
timestamp 1657128861
transform 1 0 796 0 1 600
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
timestamp 1657128861
transform 1 0 0 0 1 600
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1657128861
transform 1 0 4887 0 1 335
box 0 0 796 796
use sky130_fd_pr__res_high_po_1p41_LKUZST  XR3
timestamp 1662486269
transform 1 0 63910 0 1 100
box -307 -1408 307 1408
use sky130_fd_pr__res_high_po_1p41_S8KB58  XR4
timestamp 1662486269
transform 1 0 63349 0 1 3582
box -307 -4837 307 4837
use sky130_fd_pr__res_high_po_1p41_6AVB5Q  XR_porst
timestamp 1662486269
transform 1 0 64471 0 1 837
box -307 -2198 307 2198
use sky130_fd_pr__res_high_po_1p41_7S2UWS  XRref_high
timestamp 1662486269
transform 1 0 62788 0 1 14746
box -307 -15948 307 15948
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh1
timestamp 1662486269
transform 1 0 57520 0 1 10008
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh2
timestamp 1662486269
transform 1 0 58945 0 1 9955
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh3
timestamp 1662486269
transform 1 0 60370 0 1 9902
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh4
timestamp 1662486269
transform 1 0 61795 0 1 9849
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh
timestamp 1662486269
transform 1 0 56095 0 1 10061
box -739 -10998 739 10998
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0 ~/project/sloci/design/layout/magic_devices/opamp_layout
timestamp 1662486559
transform 1 0 26428 0 1 5058
box -5380 520 6776 6403
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_1
timestamp 1662486559
transform 1 0 26486 0 1 -1368
box -5380 520 6776 6403
<< end >>
