magic
tech sky130A
magscale 1 2
timestamp 1662393407
<< metal1 >>
rect 212 5342 222 5462
rect 302 5342 312 5462
rect 396 5449 442 5465
rect 396 4380 402 5449
rect 436 4380 442 5449
rect 528 5342 538 5462
rect 618 5342 628 5462
rect 712 5449 758 5461
rect 52 4260 62 4380
rect 142 4260 152 4380
rect 368 4260 378 4380
rect 458 4260 468 4380
rect 554 4273 560 5342
rect 594 4277 600 5342
rect 712 4380 718 5449
rect 752 4380 758 5449
rect 844 5342 854 5462
rect 934 5342 944 5462
rect 1028 5449 1074 5461
rect 568 4273 600 4277
rect 554 4261 600 4273
rect 684 4260 694 4380
rect 774 4260 784 4380
rect 870 4273 876 5342
rect 910 4273 916 5342
rect 1028 4380 1034 5449
rect 1068 4380 1074 5449
rect 1160 5342 1170 5462
rect 1250 5342 1260 5462
rect 1344 5449 1390 5465
rect 870 4261 916 4273
rect 1000 4260 1010 4380
rect 1090 4260 1100 4380
rect 1186 4273 1192 5342
rect 1226 4273 1232 5342
rect 1344 4380 1350 5449
rect 1384 4380 1390 5449
rect 1476 5342 1486 5462
rect 1566 5342 1576 5462
rect 1660 5449 1706 5461
rect 1186 4261 1232 4273
rect 1316 4260 1326 4380
rect 1406 4260 1416 4380
rect 1502 4273 1508 5342
rect 1542 4277 1548 5342
rect 1660 4380 1666 5449
rect 1700 4380 1706 5449
rect 1792 5342 1802 5462
rect 1882 5342 1892 5462
rect 1976 5449 2022 5461
rect 1516 4273 1548 4277
rect 1502 4261 1548 4273
rect 1632 4260 1642 4380
rect 1722 4260 1732 4380
rect 1818 4273 1824 5342
rect 1858 4273 1864 5342
rect 1976 4380 1982 5449
rect 2016 4380 2022 5449
rect 2108 5342 2118 5462
rect 2198 5342 2208 5462
rect 2292 5449 2338 5465
rect 1818 4261 1864 4273
rect 1948 4260 1958 4380
rect 2038 4260 2048 4380
rect 2134 4273 2140 5342
rect 2174 4273 2180 5342
rect 2292 4380 2298 5449
rect 2332 4380 2338 5449
rect 2134 4261 2180 4273
rect 2264 4260 2274 4380
rect 2354 4260 2364 4380
rect -140 4214 -70 4220
rect -140 4180 142 4214
rect -140 2850 -70 4180
rect 147 4174 2293 4220
rect 80 4085 126 4097
rect 80 3016 86 4085
rect 120 3016 126 4085
rect 212 3978 222 4098
rect 302 3978 312 4098
rect 396 4085 442 4101
rect 52 2896 62 3016
rect 142 2896 152 3016
rect 238 2909 244 3978
rect 278 2909 284 3978
rect 396 3016 402 4085
rect 436 3016 442 4085
rect 528 3978 538 4098
rect 618 3978 628 4098
rect 712 4085 758 4097
rect 238 2897 284 2909
rect 368 2896 378 3016
rect 458 2896 468 3016
rect 554 2909 560 3978
rect 594 2913 600 3978
rect 712 3016 718 4085
rect 752 3016 758 4085
rect 844 3978 854 4098
rect 934 3978 944 4098
rect 1028 4085 1074 4097
rect 568 2909 600 2913
rect 554 2897 600 2909
rect 684 2896 694 3016
rect 774 2896 784 3016
rect 870 2909 876 3978
rect 910 2909 916 3978
rect 1028 3016 1034 4085
rect 1068 3016 1074 4085
rect 1160 3978 1170 4098
rect 1250 3978 1260 4098
rect 1344 4085 1390 4101
rect 870 2897 916 2909
rect 1000 2896 1010 3016
rect 1090 2896 1100 3016
rect 1186 2909 1192 3978
rect 1226 2909 1232 3978
rect 1344 3016 1350 4085
rect 1384 3016 1390 4085
rect 1476 3978 1486 4098
rect 1566 3978 1576 4098
rect 1660 4085 1706 4097
rect 1186 2897 1232 2909
rect 1316 2896 1326 3016
rect 1406 2896 1416 3016
rect 1502 2909 1508 3978
rect 1542 2913 1548 3978
rect 1660 3016 1666 4085
rect 1700 3016 1706 4085
rect 1792 3978 1802 4098
rect 1882 3978 1892 4098
rect 1976 4085 2022 4097
rect 1516 2909 1548 2913
rect 1502 2897 1548 2909
rect 1632 2896 1642 3016
rect 1722 2896 1732 3016
rect 1818 2909 1824 3978
rect 1858 2909 1864 3978
rect 1976 3016 1982 4085
rect 2016 3016 2022 4085
rect 2108 3978 2118 4098
rect 2198 3978 2208 4098
rect 2292 4085 2338 4101
rect 1818 2897 1864 2909
rect 1948 2896 1958 3016
rect 2038 2896 2048 3016
rect 2134 2909 2140 3978
rect 2174 2909 2180 3978
rect 2292 3016 2298 4085
rect 2332 3016 2338 4085
rect 2134 2897 2180 2909
rect 2264 2896 2274 3016
rect 2354 2896 2364 3016
rect -140 2816 142 2850
rect -140 1484 -70 2816
rect 147 2809 2293 2855
rect 80 2719 126 2731
rect 80 1650 86 2719
rect 120 1650 126 2719
rect 212 2612 222 2732
rect 302 2612 312 2732
rect 396 2719 442 2735
rect 52 1530 62 1650
rect 142 1530 152 1650
rect 238 1543 244 2612
rect 278 1543 284 2612
rect 396 1650 402 2719
rect 436 1650 442 2719
rect 528 2612 538 2732
rect 618 2612 628 2732
rect 712 2719 758 2731
rect 238 1531 284 1543
rect 368 1530 378 1650
rect 458 1530 468 1650
rect 554 1543 560 2612
rect 594 1547 600 2612
rect 712 1650 718 2719
rect 752 1650 758 2719
rect 844 2612 854 2732
rect 934 2612 944 2732
rect 1028 2719 1074 2731
rect 568 1543 600 1547
rect 554 1531 600 1543
rect 684 1530 694 1650
rect 774 1530 784 1650
rect 870 1543 876 2612
rect 910 1543 916 2612
rect 1028 1650 1034 2719
rect 1068 1650 1074 2719
rect 1160 2612 1170 2732
rect 1250 2612 1260 2732
rect 1344 2719 1390 2735
rect 870 1531 916 1543
rect 1000 1530 1010 1650
rect 1090 1530 1100 1650
rect 1186 1543 1192 2612
rect 1226 1543 1232 2612
rect 1344 1650 1350 2719
rect 1384 1650 1390 2719
rect 1476 2612 1486 2732
rect 1566 2612 1576 2732
rect 1660 2719 1706 2731
rect 1186 1531 1232 1543
rect 1316 1530 1326 1650
rect 1406 1530 1416 1650
rect 1502 1543 1508 2612
rect 1542 1547 1548 2612
rect 1660 1650 1666 2719
rect 1700 1650 1706 2719
rect 1792 2612 1802 2732
rect 1882 2612 1892 2732
rect 1976 2719 2022 2731
rect 1516 1543 1548 1547
rect 1502 1531 1548 1543
rect 1632 1530 1642 1650
rect 1722 1530 1732 1650
rect 1818 1543 1824 2612
rect 1858 1543 1864 2612
rect 1976 1650 1982 2719
rect 2016 1650 2022 2719
rect 2108 2612 2118 2732
rect 2198 2612 2208 2732
rect 2292 2719 2338 2735
rect 1818 1531 1864 1543
rect 1948 1530 1958 1650
rect 2038 1530 2048 1650
rect 2134 1543 2140 2612
rect 2174 1543 2180 2612
rect 2292 1650 2298 2719
rect 2332 1650 2338 2719
rect 2134 1531 2180 1543
rect 2264 1530 2274 1650
rect 2354 1530 2364 1650
rect -140 1450 142 1484
rect -140 118 -70 1450
rect 147 1444 2293 1490
rect 80 1353 126 1365
rect 80 284 86 1353
rect 120 284 126 1353
rect 212 1246 222 1366
rect 302 1246 312 1366
rect 396 1353 442 1369
rect 52 164 62 284
rect 142 164 152 284
rect 238 177 244 1246
rect 278 177 284 1246
rect 396 284 402 1353
rect 436 284 442 1353
rect 528 1246 538 1366
rect 618 1246 628 1366
rect 712 1353 758 1365
rect 238 165 284 177
rect 368 164 378 284
rect 458 164 468 284
rect 554 177 560 1246
rect 594 181 600 1246
rect 712 284 718 1353
rect 752 284 758 1353
rect 844 1246 854 1366
rect 934 1246 944 1366
rect 1028 1353 1074 1365
rect 568 177 600 181
rect 554 165 600 177
rect 684 164 694 284
rect 774 164 784 284
rect 870 177 876 1246
rect 910 177 916 1246
rect 1028 284 1034 1353
rect 1068 284 1074 1353
rect 1160 1246 1170 1366
rect 1250 1246 1260 1366
rect 1344 1353 1390 1369
rect 870 165 916 177
rect 1000 164 1010 284
rect 1090 164 1100 284
rect 1186 177 1192 1246
rect 1226 177 1232 1246
rect 1344 284 1350 1353
rect 1384 284 1390 1353
rect 1476 1246 1486 1366
rect 1566 1246 1576 1366
rect 1660 1353 1706 1365
rect 1186 165 1232 177
rect 1316 164 1326 284
rect 1406 164 1416 284
rect 1502 177 1508 1246
rect 1542 181 1548 1246
rect 1660 284 1666 1353
rect 1700 284 1706 1353
rect 1792 1246 1802 1366
rect 1882 1246 1892 1366
rect 1976 1353 2022 1365
rect 1516 177 1548 181
rect 1502 165 1548 177
rect 1632 164 1642 284
rect 1722 164 1732 284
rect 1818 177 1824 1246
rect 1858 177 1864 1246
rect 1976 284 1982 1353
rect 2016 284 2022 1353
rect 2108 1246 2118 1366
rect 2198 1246 2208 1366
rect 2292 1353 2338 1369
rect 1818 165 1864 177
rect 1948 164 1958 284
rect 2038 164 2048 284
rect 2134 177 2140 1246
rect 2174 177 2180 1246
rect 2292 284 2298 1353
rect 2332 284 2338 1353
rect 2134 165 2180 177
rect 2264 164 2274 284
rect 2354 164 2364 284
rect -140 84 142 118
rect -140 80 -70 84
rect 147 79 2293 125
<< via1 >>
rect 222 5342 302 5462
rect 538 5342 618 5462
rect 62 4260 142 4380
rect 378 4260 458 4380
rect 854 5342 934 5462
rect 694 4260 774 4380
rect 1170 5342 1250 5462
rect 1010 4260 1090 4380
rect 1486 5342 1566 5462
rect 1326 4260 1406 4380
rect 1802 5342 1882 5462
rect 1642 4260 1722 4380
rect 2118 5342 2198 5462
rect 1958 4260 2038 4380
rect 2274 4260 2354 4380
rect 222 3978 302 4098
rect 62 2896 142 3016
rect 538 3978 618 4098
rect 378 2896 458 3016
rect 854 3978 934 4098
rect 694 2896 774 3016
rect 1170 3978 1250 4098
rect 1010 2896 1090 3016
rect 1486 3978 1566 4098
rect 1326 2896 1406 3016
rect 1802 3978 1882 4098
rect 1642 2896 1722 3016
rect 2118 3978 2198 4098
rect 1958 2896 2038 3016
rect 2274 2896 2354 3016
rect 222 2612 302 2732
rect 62 1530 142 1650
rect 538 2612 618 2732
rect 378 1530 458 1650
rect 854 2612 934 2732
rect 694 1530 774 1650
rect 1170 2612 1250 2732
rect 1010 1530 1090 1650
rect 1486 2612 1566 2732
rect 1326 1530 1406 1650
rect 1802 2612 1882 2732
rect 1642 1530 1722 1650
rect 2118 2612 2198 2732
rect 1958 1530 2038 1650
rect 2274 1530 2354 1650
rect 222 1246 302 1366
rect 62 164 142 284
rect 538 1246 618 1366
rect 378 164 458 284
rect 854 1246 934 1366
rect 694 164 774 284
rect 1170 1246 1250 1366
rect 1010 164 1090 284
rect 1486 1246 1566 1366
rect 1326 164 1406 284
rect 1802 1246 1882 1366
rect 1642 164 1722 284
rect 2118 1246 2198 1366
rect 1958 164 2038 284
rect 2274 164 2354 284
<< metal2 >>
rect 222 5462 2198 5472
rect 302 5342 538 5462
rect 618 5342 854 5462
rect 934 5460 1170 5462
rect 1250 5460 1486 5462
rect 934 5360 1140 5460
rect 1280 5360 1486 5460
rect 934 5342 1170 5360
rect 1250 5342 1486 5360
rect 1566 5342 1802 5462
rect 1882 5342 2118 5462
rect 222 5332 2198 5342
rect -40 4380 2354 4390
rect -40 4260 62 4380
rect 142 4260 378 4380
rect 458 4260 694 4380
rect 774 4260 1010 4380
rect 1090 4260 1326 4380
rect 1406 4260 1642 4380
rect 1722 4260 1958 4380
rect 2038 4260 2274 4380
rect -40 4250 2354 4260
rect -40 3026 140 4250
rect 222 4098 2198 4108
rect 302 3978 538 4098
rect 618 3978 854 4098
rect 934 4080 1170 4098
rect 1250 4080 1486 4098
rect 934 3980 1140 4080
rect 1280 3980 1486 4080
rect 934 3978 1170 3980
rect 1250 3978 1486 3980
rect 1566 3978 1802 4098
rect 1882 3978 2118 4098
rect 222 3968 2198 3978
rect -40 3016 2354 3026
rect -40 2896 62 3016
rect 142 2896 378 3016
rect 458 2896 694 3016
rect 774 2896 1010 3016
rect 1090 2896 1326 3016
rect 1406 2896 1642 3016
rect 1722 2896 1958 3016
rect 2038 2896 2274 3016
rect -40 2886 2354 2896
rect -40 1660 140 2886
rect 222 2732 2198 2742
rect 302 2612 538 2732
rect 618 2612 854 2732
rect 934 2720 1170 2732
rect 1250 2720 1486 2732
rect 934 2620 1140 2720
rect 1280 2620 1486 2720
rect 934 2612 1170 2620
rect 1250 2612 1486 2620
rect 1566 2612 1802 2732
rect 1882 2612 2118 2732
rect 222 2602 2198 2612
rect -40 1650 2354 1660
rect -40 1530 62 1650
rect 142 1530 378 1650
rect 458 1530 694 1650
rect 774 1530 1010 1650
rect 1090 1530 1326 1650
rect 1406 1530 1642 1650
rect 1722 1530 1958 1650
rect 2038 1530 2274 1650
rect -40 1520 2354 1530
rect -40 294 140 1520
rect 222 1366 2198 1376
rect 302 1246 538 1366
rect 618 1246 854 1366
rect 934 1360 1170 1366
rect 1250 1360 1486 1366
rect 934 1246 1140 1360
rect 1280 1246 1486 1360
rect 1566 1246 1802 1366
rect 1882 1246 2118 1366
rect 222 1240 1140 1246
rect 1280 1240 2198 1246
rect 222 1236 2198 1240
rect 1140 1230 1280 1236
rect -40 284 2354 294
rect -40 164 62 284
rect 142 164 378 284
rect 458 164 694 284
rect 774 164 1010 284
rect 1090 164 1326 284
rect 1406 164 1642 284
rect 1722 164 1958 284
rect 2038 164 2274 284
rect -40 154 2354 164
rect -40 150 140 154
<< via2 >>
rect 1140 5360 1170 5460
rect 1170 5360 1250 5460
rect 1250 5360 1280 5460
rect 1140 3980 1170 4080
rect 1170 3980 1250 4080
rect 1250 3980 1280 4080
rect 1140 2620 1170 2720
rect 1170 2620 1250 2720
rect 1250 2620 1280 2720
rect 1140 1246 1170 1360
rect 1170 1246 1250 1360
rect 1250 1246 1280 1360
rect 1140 1240 1280 1246
<< metal3 >>
rect 1130 5460 1290 5650
rect 1130 5360 1140 5460
rect 1280 5360 1290 5460
rect 1130 4080 1290 5360
rect 1130 3980 1140 4080
rect 1280 3980 1290 4080
rect 1130 2720 1290 3980
rect 1130 2620 1140 2720
rect 1280 2620 1290 2720
rect 1130 1360 1290 2620
rect 1130 1240 1140 1360
rect 1280 1240 1290 1360
rect 1130 1235 1290 1240
use sky130_fd_pr__pfet_01v8_lvt_D74VRS  sky130_fd_pr__pfet_01v8_lvt_D74VRS_0
timestamp 1661879915
transform 1 0 1209 0 1 2778
box -1273 -2831 1273 2831
<< end >>
