magic
tech sky130A
magscale 1 2
timestamp 1661906430
<< metal1 >>
rect 517 1023 527 1113
rect 617 1023 627 1113
rect 1007 1101 1053 1113
rect 1007 801 1013 1101
rect 1047 801 1053 1101
rect 1433 1023 1443 1113
rect 1533 1023 1543 1113
rect 1923 1101 1969 1113
rect 59 711 69 801
rect 159 711 169 801
rect 975 711 985 801
rect 1075 711 1085 801
rect 1465 725 1471 1023
rect 1505 725 1511 1023
rect 1923 801 1929 1101
rect 1963 801 1969 1101
rect 2349 1023 2359 1113
rect 2449 1023 2459 1113
rect 1465 713 1511 725
rect 1891 711 1901 801
rect 1991 711 2001 801
rect 2381 725 2387 1023
rect 2421 725 2427 1023
rect 2381 713 2427 725
rect 527 635 617 681
rect 985 635 1075 681
rect 1443 635 1533 681
rect 1901 635 1991 681
rect 91 545 137 557
rect 91 245 97 545
rect 131 245 137 545
rect 517 467 527 557
rect 617 467 627 557
rect 1007 545 1053 557
rect 59 155 69 245
rect 159 155 169 245
rect 549 169 555 467
rect 589 169 595 467
rect 1007 245 1013 545
rect 1047 245 1053 545
rect 1433 467 1443 557
rect 1533 467 1543 557
rect 1923 545 1969 557
rect 549 157 595 169
rect 975 155 985 245
rect 1075 155 1085 245
rect 1465 169 1471 467
rect 1505 169 1511 467
rect 1923 245 1929 545
rect 1963 245 1969 545
rect 2349 467 2359 557
rect 2449 467 2459 557
rect 1465 157 1511 169
rect 1891 155 1901 245
rect 1991 155 2001 245
rect 2381 169 2387 467
rect 2421 169 2427 467
rect 2381 157 2427 169
rect 527 79 617 125
rect 985 79 1075 125
rect 1443 79 1533 125
rect 1901 79 1991 125
<< via1 >>
rect 527 1023 617 1113
rect 1443 1023 1533 1113
rect 69 711 159 801
rect 985 711 1075 801
rect 2359 1023 2449 1113
rect 1901 711 1991 801
rect 527 467 617 557
rect 69 155 159 245
rect 1443 467 1533 557
rect 985 155 1075 245
rect 2359 467 2449 557
rect 1901 155 1991 245
<< metal2 >>
rect 527 1113 2449 1123
rect 617 1023 1443 1113
rect 1533 1023 2359 1113
rect 527 1013 2449 1023
rect 69 801 1991 811
rect 159 711 985 801
rect 1075 711 1901 801
rect 69 701 1991 711
rect 527 557 617 567
rect 527 457 617 467
rect 1443 557 1533 567
rect 1443 457 1533 467
rect 2359 557 2449 567
rect 2359 457 2449 467
rect 69 245 159 255
rect 69 145 159 155
rect 985 245 1075 255
rect 985 145 1075 155
rect 1901 245 1991 255
rect 1901 145 1991 155
use sky130_fd_pr__nfet_01v8_lvt_UV2JYN  sky130_fd_pr__nfet_01v8_lvt_UV2JYN_0
timestamp 1661905147
transform 1 0 1259 0 1 604
box -1312 -657 1312 657
<< end >>
