magic
tech sky130A
magscale 1 2
timestamp 1662733787
use sky130_fd_pr__cap_mim_m3_1_Y9W37A  sky130_fd_pr__cap_mim_m3_1_Y9W37A_0
timestamp 1662733733
transform 1 0 3182 0 1 526
box -2450 -680 2318 680
use sky130_fd_pr__nfet_01v8_Y5UG24  sky130_fd_pr__nfet_01v8_Y5UG24_0
timestamp 1662731509
transform 1 0 194 0 1 -387
box -246 -329 246 329
use sky130_fd_pr__nfet_01v8_Y5UG24  sky130_fd_pr__nfet_01v8_Y5UG24_1
timestamp 1662731509
transform 1 0 580 0 1 -387
box -246 -329 246 329
use sky130_fd_pr__nfet_01v8_Y5UG24  sky130_fd_pr__nfet_01v8_Y5UG24_2
timestamp 1662731509
transform 1 0 966 0 1 -387
box -246 -329 246 329
use sky130_fd_pr__pfet_01v8_TSNZVH  sky130_fd_pr__pfet_01v8_TSNZVH_0
timestamp 1662731045
transform 1 0 193 0 1 531
box -246 -584 246 584
use sky130_fd_pr__pfet_01v8_TSNZVH  sky130_fd_pr__pfet_01v8_TSNZVH_1
timestamp 1662731045
transform 1 0 580 0 1 532
box -246 -584 246 584
use sky130_fd_pr__res_high_po_1p41_2TBR6S  sky130_fd_pr__res_high_po_1p41_2TBR6S_0
timestamp 1662731843
transform 0 1 3304 -1 0 -411
box -307 -2198 307 2198
<< end >>
