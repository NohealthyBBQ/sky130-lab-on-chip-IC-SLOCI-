magic
tech sky130A
magscale 1 2
timestamp 1661881632
<< metal1 >>
rect 212 5342 222 5462
rect 302 5342 312 5462
rect 396 5453 442 5465
rect 396 4384 402 5453
rect 436 4384 442 5453
rect 528 5346 538 5466
rect 618 5346 628 5466
rect 52 4260 62 4380
rect 142 4260 152 4380
rect 368 4264 378 4384
rect 458 4264 468 4384
rect 554 4277 560 5346
rect 594 4277 600 5346
rect 554 4265 600 4277
rect 147 4174 2293 4220
rect 147 2809 2293 2855
rect 147 1444 2293 1490
rect 147 79 2293 125
<< via1 >>
rect 222 5342 302 5462
rect 538 5346 618 5466
rect 62 4260 142 4380
rect 378 4264 458 4384
<< metal2 >>
rect 222 5462 302 5472
rect 222 5332 302 5342
rect 538 5466 618 5476
rect 538 5336 618 5346
rect 62 4380 142 4390
rect 62 4250 142 4260
rect 378 4384 458 4394
rect 378 4254 458 4264
use sky130_fd_pr__pfet_01v8_lvt_D74VRS  sky130_fd_pr__pfet_01v8_lvt_D74VRS_0
timestamp 1661879915
transform 1 0 1209 0 1 2778
box -1273 -2831 1273 2831
<< end >>
