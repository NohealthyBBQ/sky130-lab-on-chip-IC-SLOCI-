magic
tech sky130A
magscale 1 2
timestamp 1662233295
<< metal2 >>
rect -3780 2660 -3710 2670
rect -3780 2590 -3710 2600
rect -2480 2660 -1640 2670
rect -2480 2600 -1740 2660
rect -1670 2600 -1640 2660
rect -2480 2590 -1640 2600
<< via2 >>
rect -3780 2600 -3710 2660
rect -1740 2600 -1670 2660
<< metal3 >>
rect -3832 2665 -3702 4230
rect -3832 2660 -3700 2665
rect -3832 2600 -3780 2660
rect -3710 2600 -3700 2660
rect -3832 2595 -3700 2600
rect -1772 2660 -1642 4038
rect -1772 2600 -1740 2660
rect -1670 2600 -1642 2660
rect -3832 2590 -3702 2595
rect -1772 2560 -1642 2600
use XM_actload2  XM_actload2_0
timestamp 1661870098
transform 1 0 2789 0 1 -857
box -53 -53 2571 3173
use XM_cs  XM_cs_0
timestamp 1661891635
transform 1 0 6296 0 1 3675
box -64 -53 2482 5609
use XM_diffpair  XM_diffpair_0
timestamp 1662136735
transform 1 0 -3688 0 1 2162
box -400 -1642 1600 1820
use XM_ppair  XM_ppair_0
timestamp 1662231221
transform 1 0 -5102 0 1 5030
box -220 -1160 4440 828
use XM_tail  XM_tail_0
timestamp 1661906530
transform 1 0 615 0 1 4879
box -53 -53 2571 1261
use sky130_fd_pr__cap_mim_m3_1_EN3Q86  sky130_fd_pr__cap_mim_m3_1_EN3Q86_0
timestamp 1661639644
transform 1 0 8170 0 1 724
box -1750 -2240 1749 2240
use sky130_fd_pr__res_high_po_2p85_7J2RPB  sky130_fd_pr__res_high_po_2p85_7J2RPB_0
timestamp 1662230297
transform 1 0 12090 0 1 4991
box -451 -1808 451 1808
<< end >>
