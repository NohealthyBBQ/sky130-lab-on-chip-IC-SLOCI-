magic
tech sky130A
magscale 1 2
timestamp 1662719632
<< nwell >>
rect -140 -160 2080 1600
<< nsubdiff >>
rect -60 1520 2000 1560
rect -60 -80 2000 -40
<< locali >>
rect -60 1520 2000 1560
rect -60 -80 2000 -40
<< metal1 >>
rect 30 1340 40 1400
rect 100 1340 110 1400
rect 550 1340 560 1400
rect 620 1340 630 1400
rect 1070 1340 1080 1400
rect 1140 1340 1150 1400
rect 1570 1340 1580 1400
rect 1640 1340 1650 1400
rect 290 1200 300 1260
rect 360 1200 370 1260
rect 810 1200 820 1260
rect 880 1200 890 1260
rect 1330 1200 1340 1260
rect 1400 1200 1410 1260
rect 1830 1200 1840 1260
rect 1900 1200 1910 1260
rect 104 1108 1842 1154
rect 30 980 40 1040
rect 100 980 110 1040
rect 550 980 560 1040
rect 620 980 630 1040
rect 1070 980 1080 1040
rect 1140 980 1150 1040
rect 1570 980 1580 1040
rect 1640 980 1650 1040
rect 290 820 300 880
rect 360 820 370 880
rect 810 820 820 880
rect 880 820 890 880
rect 1310 820 1320 880
rect 1380 820 1390 880
rect 1830 820 1840 880
rect 1900 820 1910 880
rect 102 742 1840 788
rect 30 600 40 660
rect 100 600 110 660
rect 550 600 560 660
rect 620 600 630 660
rect 1050 600 1060 660
rect 1120 600 1130 660
rect 1570 600 1580 660
rect 1640 600 1650 660
rect 290 460 300 520
rect 360 460 370 520
rect 790 460 800 520
rect 860 460 870 520
rect 1310 460 1320 520
rect 1380 460 1390 520
rect 1830 460 1840 520
rect 1900 460 1910 520
rect 100 382 1838 428
rect 30 240 40 300
rect 100 240 110 300
rect 550 240 560 300
rect 620 240 630 300
rect 1050 240 1060 300
rect 1120 240 1130 300
rect 1570 240 1580 300
rect 1640 240 1650 300
rect 290 100 300 160
rect 360 100 370 160
rect 790 100 800 160
rect 860 100 870 160
rect 1310 100 1320 160
rect 1380 100 1390 160
rect 1830 100 1840 160
rect 1900 100 1910 160
rect 102 14 1840 60
<< via1 >>
rect 40 1340 100 1400
rect 560 1340 620 1400
rect 1080 1340 1140 1400
rect 1580 1340 1640 1400
rect 300 1200 360 1260
rect 820 1200 880 1260
rect 1340 1200 1400 1260
rect 1840 1200 1900 1260
rect 40 980 100 1040
rect 560 980 620 1040
rect 1080 980 1140 1040
rect 1580 980 1640 1040
rect 300 820 360 880
rect 820 820 880 880
rect 1320 820 1380 880
rect 1840 820 1900 880
rect 40 600 100 660
rect 560 600 620 660
rect 1060 600 1120 660
rect 1580 600 1640 660
rect 300 460 360 520
rect 800 460 860 520
rect 1320 460 1380 520
rect 1840 460 1900 520
rect 40 240 100 300
rect 560 240 620 300
rect 1060 240 1120 300
rect 1580 240 1640 300
rect 300 100 360 160
rect 800 100 860 160
rect 1320 100 1380 160
rect 1840 100 1900 160
<< metal2 >>
rect 40 1400 100 1410
rect 560 1400 620 1410
rect 1080 1400 1140 1410
rect 1580 1400 1640 1410
rect 100 1340 560 1400
rect 620 1340 1080 1400
rect 1140 1340 1580 1400
rect 40 1040 100 1340
rect 560 1330 620 1340
rect 1080 1330 1140 1340
rect 1580 1330 1640 1340
rect 300 1260 360 1270
rect 820 1260 880 1270
rect 1340 1260 1400 1270
rect 1840 1260 1900 1270
rect 360 1200 820 1260
rect 880 1200 1340 1260
rect 1400 1200 1840 1260
rect 300 1190 360 1200
rect 820 1190 880 1200
rect 1340 1190 1400 1200
rect 560 1040 620 1050
rect 1080 1040 1140 1050
rect 1580 1040 1640 1050
rect 100 980 560 1040
rect 620 980 1080 1040
rect 1140 980 1580 1040
rect 40 660 100 980
rect 560 970 620 980
rect 1080 970 1140 980
rect 1580 970 1640 980
rect 300 880 360 890
rect 820 880 880 890
rect 1320 880 1380 890
rect 1840 880 1900 1200
rect 360 820 820 880
rect 880 820 1320 880
rect 1380 820 1840 880
rect 300 810 360 820
rect 820 810 880 820
rect 1320 810 1380 820
rect 560 660 620 670
rect 1060 660 1120 670
rect 1580 660 1640 670
rect 100 600 560 660
rect 620 600 1060 660
rect 1120 600 1580 660
rect 40 300 100 600
rect 560 590 620 600
rect 1060 590 1120 600
rect 1580 590 1640 600
rect 300 520 360 530
rect 800 520 860 530
rect 1320 520 1380 530
rect 1840 520 1900 820
rect 360 460 800 520
rect 860 460 1320 520
rect 1380 460 1840 520
rect 300 450 360 460
rect 800 450 860 460
rect 1320 450 1380 460
rect 560 300 620 310
rect 1060 300 1120 310
rect 1580 300 1640 310
rect 100 240 560 300
rect 620 240 1060 300
rect 1120 240 1580 300
rect 40 230 100 240
rect 560 230 620 240
rect 1060 230 1120 240
rect 1580 230 1640 240
rect 300 160 360 170
rect 800 160 860 170
rect 1320 160 1380 170
rect 1840 160 1900 460
rect 360 100 800 160
rect 860 100 1320 160
rect 1380 100 1840 160
rect 300 90 360 100
rect 800 90 860 100
rect 1320 90 1380 100
rect 1840 90 1900 100
use sky130_fd_pr__pfet_01v8_lvt_9UM225  sky130_fd_pr__pfet_01v8_lvt_9UM225_0
timestamp 1662718844
transform 1 0 968 0 1 712
box -968 -712 968 745
<< end >>
