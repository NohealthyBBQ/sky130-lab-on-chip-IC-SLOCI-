** sch_path: /foss/designs/sumprj/hiarachy_final/buffer_amp_vop.sch
.subckt buffer_amp_vop BIAS GND SUB I1A I1B I2A I2B I3A I3B I4A I4B VDD AMP VOP OUT0 OUT180 OUT90
+ OUT270
*.PININFO BIAS:I GND:I SUB:I I1A:I I1B:I I2A:I I2B:I I3A:I I3B:I I4A:I I4B:I VDD:I AMP:O VOP:O
*+ OUT0:O OUT180:O OUT90:O OUT270:O
X2 I2A I2B BIAS VDD GND SUB net1 net1 buffer_amp
X4 I4A I4B BIAS VDD GND SUB net1 net1 buffer_amp
X1 I1A I1B BIAS VDD GND SUB OUT0 OUT180 buffer_amp
X3 I3A I3B BIAS VDD GND SUB OUT90 OUT270 buffer_amp
X5 OUT180 OUT0 OUT90 OUT270 AMP VDD GND SUB amp_dec
X6 net1 VDD GND SUB VOP vop_dec
.ends

* expanding   symbol:  hiarachy_final/buffer_amp.sym # of pins=8
** sym_path: /foss/designs/sumprj/hiarachy_final/buffer_amp.sym
** sch_path: /foss/designs/sumprj/hiarachy_final/buffer_amp.sch
.subckt buffer_amp  INA INB BIAS VDD GND SUB OUTA OUTB
*.PININFO INA:I INB:I BIAS:I GND:I VDD:I SUB:I OUTA:O OUTB:O
XM1 net1 BIAS GND SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUTB INB net1 SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUTA INA net1 SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR2 OUTB VDD SUB sky130_fd_pr__res_high_po_5p73 L=30.4 mult=1 m=1
XR1 OUTA VDD SUB sky130_fd_pr__res_high_po_5p73 L=30.4 mult=1 m=1
XM4 net1 BIAS GND SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  hiarachy_final/amp_dec.sym # of pins=8
** sym_path: /foss/designs/sumprj/hiarachy_final/amp_dec.sym
** sch_path: /foss/designs/sumprj/hiarachy_final/amp_dec.sch
.subckt amp_dec  IN1 IN2 IN3 IN4 AMP VDD GND SUB
*.PININFO VDD:I SUB:I GND:I IN1:I IN2:I IN3:I IN4:I AMP:O
XM25 VDD IN1 AMP SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 AMP GND sky130_fd_pr__cap_mim_m3_1 W=20 L=30 MF=1 m=1
XM26 VDD IN2 AMP SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM27 VDD IN3 AMP SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM28 VDD IN4 AMP SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR18 GND AMP SUB sky130_fd_pr__res_high_po_2p85 L=42 mult=1 m=1
.ends


* expanding   symbol:  hiarachy_final/vop_dec.sym # of pins=5
** sym_path: /foss/designs/sumprj/hiarachy_final/vop_dec.sym
** sch_path: /foss/designs/sumprj/hiarachy_final/vop_dec.sch
.subckt vop_dec  IN VDD GND SUB VOP
*.PININFO IN:I VDD:I GND:I SUB:I VOP:O
XM41 VDD IN VOP SUB sky130_fd_pr__nfet_01v8_lvt L=0.15 W=12 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC2 IN GND sky130_fd_pr__cap_mim_m3_1 W=20 L=30 MF=1 m=1
XR21 GND VOP SUB sky130_fd_pr__res_high_po_2p85 L=42 mult=1 m=1
.ends

.end
