magic
tech sky130A
magscale 1 2
timestamp 1662515827
<< locali >>
rect 6430 9730 6730 9770
rect 6430 8350 6730 8390
<< metal1 >>
rect 5770 9810 6340 9830
rect 5770 9420 5780 9810
rect 6320 9420 6340 9810
rect 5770 9400 6340 9420
rect 6780 8400 6840 9670
rect 6870 9610 7000 9670
rect 7060 9610 7070 9670
rect 6990 9600 7070 9610
rect 6870 9510 6880 9570
rect 6940 9520 7070 9570
rect 6940 9510 6950 9520
rect 6870 9500 6950 9510
rect 6990 9470 7000 9480
rect 6870 9420 7000 9470
rect 7060 9420 7070 9480
rect 6990 9410 7070 9420
rect 6870 9320 6880 9380
rect 6940 9320 7070 9380
rect 6870 9310 6950 9320
rect 6990 9280 7000 9290
rect 6870 9230 7000 9280
rect 7060 9230 7070 9290
rect 6990 9220 7070 9230
rect 6870 9130 6880 9190
rect 6940 9180 6950 9190
rect 6940 9130 7070 9180
rect 6870 9120 6950 9130
rect 6870 9040 7000 9090
rect 6990 9030 7000 9040
rect 7060 9030 7070 9090
rect 6990 9020 7070 9030
rect 6870 8940 6880 9000
rect 6940 8990 6950 9000
rect 6940 8940 7070 8990
rect 6870 8930 6950 8940
rect 6870 8850 7000 8900
rect 6990 8840 7000 8850
rect 7060 8840 7070 8900
rect 6990 8830 7070 8840
rect 6870 8750 6880 8810
rect 6940 8800 6950 8810
rect 6940 8750 7070 8800
rect 6870 8740 6950 8750
rect 6990 8700 7000 8710
rect 6870 8650 7000 8700
rect 7060 8650 7070 8710
rect 6990 8640 7070 8650
rect 6870 8550 6880 8610
rect 6940 8560 7070 8610
rect 6940 8550 6950 8560
rect 6870 8540 6950 8550
rect 6870 8460 7000 8510
rect 6990 8450 7000 8460
rect 7060 8450 7070 8510
rect 6990 8440 7070 8450
rect 7100 8400 7160 9680
rect 7420 8410 7860 8420
rect 7420 8400 7440 8410
rect 6780 8340 7440 8400
rect 7420 8320 7440 8340
rect 7840 8320 7860 8410
rect 7420 8310 7860 8320
rect 5720 1000 6380 1040
rect 5720 560 5760 1000
rect 6340 560 6380 1000
rect 5720 520 6380 560
<< via1 >>
rect 5780 9420 6320 9810
rect 7000 9610 7060 9670
rect 6880 9510 6940 9570
rect 7000 9420 7060 9480
rect 6880 9320 6940 9380
rect 7000 9230 7060 9290
rect 6880 9130 6940 9190
rect 7000 9030 7060 9090
rect 6880 8940 6940 9000
rect 7000 8840 7060 8900
rect 6880 8750 6940 8810
rect 7000 8650 7060 8710
rect 6880 8550 6940 8610
rect 7000 8450 7060 8510
rect 7440 8320 7840 8410
rect 5760 560 6340 1000
<< metal2 >>
rect 5600 9810 6950 9830
rect 5600 9420 5780 9810
rect 6320 9570 6950 9810
rect 6320 9510 6880 9570
rect 6940 9510 6950 9570
rect 6320 9420 6950 9510
rect 5600 9400 6950 9420
rect 6650 9380 6950 9400
rect 6650 9320 6880 9380
rect 6940 9320 6950 9380
rect 6650 9190 6950 9320
rect 6650 9130 6880 9190
rect 6940 9130 6950 9190
rect 6650 9000 6950 9130
rect 6650 8940 6880 9000
rect 6940 8940 6950 9000
rect 6650 8810 6950 8940
rect 6650 8750 6880 8810
rect 6940 8750 6950 8810
rect 6650 8610 6950 8750
rect 6650 8550 6880 8610
rect 6940 8550 6950 8610
rect 6650 8430 6950 8550
rect 6990 9670 7280 9990
rect 6990 9610 7000 9670
rect 7060 9610 7280 9670
rect 6990 9480 7280 9610
rect 6990 9420 7000 9480
rect 7060 9420 7280 9480
rect 6990 9290 7280 9420
rect 6990 9230 7000 9290
rect 7060 9230 7280 9290
rect 6990 9090 7280 9230
rect 6990 9030 7000 9090
rect 7060 9030 7280 9090
rect 6990 8900 7280 9030
rect 6990 8840 7000 8900
rect 7060 8840 7280 8900
rect 6990 8710 7280 8840
rect 6990 8650 7000 8710
rect 7060 8650 7280 8710
rect 6990 8510 7280 8650
rect 6990 8450 7000 8510
rect 7060 8450 7280 8510
rect 6990 8430 7280 8450
rect 7420 8410 7860 8420
rect 7420 8320 7440 8410
rect 7840 8320 7860 8410
rect 7420 8310 7860 8320
rect 5600 1000 6380 1040
rect 5600 560 5760 1000
rect 6340 560 6380 1000
rect 5600 400 6380 560
<< via2 >>
rect 7460 8320 7820 8410
rect 5760 560 6340 1000
<< metal3 >>
rect 7440 8410 7840 9990
rect 7440 8320 7460 8410
rect 7820 8320 7840 8410
rect 7440 6920 7840 8320
rect 7440 6760 7460 6920
rect 7820 6760 7840 6920
rect 7440 6740 7840 6760
rect 5720 1000 6660 1040
rect 5720 560 5760 1000
rect 6340 560 6660 1000
rect 5720 520 6660 560
<< via3 >>
rect 7460 6760 7820 6920
<< metal4 >>
rect 7440 6920 7840 6940
rect 7440 6760 7460 6920
rect 7820 6760 7840 6920
rect 7440 6080 7840 6760
use sky130_fd_pr__cap_mim_m3_1_4RCNTW  XC2 backup/1.7_10G
timestamp 1662404926
transform 1 0 8750 0 1 3500
box -2150 -3100 2149 3100
use sky130_fd_pr__nfet_01v8_lvt_6BNFGK  XM41 backup/1.7_10G
timestamp 1662404926
transform 0 1 6970 -1 0 9063
box -743 -310 743 310
use sky130_fd_pr__res_high_po_2p85_MXEQGY  XR21 backup/1.7_10G
timestamp 1662404926
transform 1 0 6051 0 1 5198
box -451 -4798 451 4798
<< labels >>
rlabel metal2 5600 400 5760 1040 1 GND
rlabel metal2 5600 9400 5780 9830 1 VOP
rlabel metal2 6990 9680 7280 9990 1 VDD
rlabel metal3 7440 8410 7840 9990 1 IN
rlabel locali 6430 8350 6730 8390 1 SUB
<< end >>
