magic
tech sky130A
magscale 1 2
timestamp 1662840447
<< nwell >>
rect -8726 10225 -8100 11452
<< locali >>
rect -1960 10600 1560 10940
rect -7740 8580 -7620 8860
rect -9000 8140 -8880 8440
rect -1960 6380 -1860 6900
rect -760 6300 -560 6900
rect 520 6320 720 6920
rect 1820 6320 2000 6920
rect 3100 6320 3300 6920
rect 4380 6320 4480 6920
<< metal1 >>
rect -7750 11040 -7740 11120
rect -7680 11040 -7670 11120
rect 1190 11100 1200 11200
rect 1300 11100 1310 11200
rect -11458 9858 -10653 9906
rect -10600 8810 -10540 11000
rect -8850 8810 -8840 8820
rect -13422 8764 -8840 8810
rect -10600 8760 -10540 8764
rect -8850 8760 -8840 8764
rect -8780 8760 -8770 8820
rect -7950 8760 -7940 8820
rect -7880 8760 -7870 8820
rect -10090 8240 -10080 8300
rect -10020 8240 -10010 8300
rect -8700 8200 -4700 8400
rect -10080 7780 -9980 7920
rect -9180 4980 -9120 7840
rect -8710 6000 -8700 6100
rect -8600 6000 -8590 6100
rect -4900 4000 -4700 8200
rect -4900 3800 -600 4000
<< via1 >>
rect -7740 11040 -7680 11120
rect 1200 11100 1300 11200
rect -8840 8760 -8780 8820
rect -7940 8760 -7880 8820
rect -10080 8240 -10020 8300
rect -8700 6000 -8600 6100
<< metal2 >>
rect 1200 11200 1300 11210
rect -8940 11120 -7680 11140
rect -8940 11040 -7740 11120
rect -8940 11020 -7680 11040
rect -14160 8460 -13540 8520
rect -14160 5760 -14100 8460
rect -11260 7680 -11180 8700
rect -10080 8300 -10020 9160
rect -8860 8840 -8760 8850
rect -8860 8730 -8760 8740
rect -8216 8840 -8114 8940
rect -8216 8820 -7880 8840
rect -8216 8760 -8200 8820
rect -8140 8760 -7940 8820
rect -8216 8740 -7880 8760
rect -10080 8230 -10020 8240
rect -11260 7620 -9480 7680
rect -9540 6100 -9480 7620
rect -8216 6980 -8114 8740
rect 1200 8700 1300 11100
rect -8700 6100 -8600 6110
rect -9540 6000 -8700 6100
rect -11600 5760 -11540 5770
rect -14160 5700 -11600 5760
rect -11600 5690 -11540 5700
rect -11460 5760 -11400 5770
rect -9540 5760 -9480 6000
rect -8700 5990 -8600 6000
rect -11400 5700 -9480 5760
rect -11460 5690 -11400 5700
rect -11460 5120 -11400 5130
rect -11460 4280 -11400 5060
rect -11520 4240 -11400 4280
rect -11620 4100 -11500 4126
rect -11620 4040 -11600 4100
rect -11540 4040 -11500 4100
rect -11620 4000 -11500 4040
rect -11280 3180 -11220 3190
rect -11280 2500 -11220 3120
rect -14220 2430 -14130 2464
rect -11280 2300 1400 2500
rect 1140 1860 1400 2300
<< via2 >>
rect -8860 8820 -8760 8840
rect -8860 8760 -8840 8820
rect -8840 8760 -8780 8820
rect -8780 8760 -8760 8820
rect -8860 8740 -8760 8760
rect -8200 8760 -8140 8820
rect -11600 5700 -11540 5760
rect -11460 5700 -11400 5760
rect -11460 5060 -11400 5120
rect -11600 4040 -11540 4100
rect -11280 3120 -11220 3180
<< metal3 >>
rect -8870 8840 -8750 8845
rect -8870 8740 -8860 8840
rect -8760 8820 -8120 8840
rect -8760 8760 -8200 8820
rect -8140 8760 -8120 8820
rect -8760 8740 -8120 8760
rect -8870 8735 -8750 8740
rect -11610 5760 -11530 5790
rect -11610 5700 -11600 5760
rect -11540 5700 -11530 5760
rect -11610 4100 -11530 5700
rect -11470 5760 -11390 5770
rect -11470 5700 -11460 5760
rect -11400 5700 -11390 5760
rect -11470 5120 -11390 5700
rect -11470 5060 -11460 5120
rect -11400 5060 -11390 5120
rect -11470 5050 -11390 5060
rect -11610 4040 -11600 4100
rect -11540 4040 -11530 4100
rect -11610 3200 -11530 4040
rect -11610 3180 -11200 3200
rect -11610 3120 -11280 3180
rect -11220 3120 -11200 3180
rect -11290 3115 -11210 3120
use XM_Rref  XM_Rref_0
timestamp 1662826901
transform 0 1 -13057 -1 0 -5305
box -1417 -1173 5029 21223
use XM_bjt  XM_bjt_0
timestamp 1662737136
transform 1 0 -1980 0 1 -2620
box 0 0 6492 9068
use XM_bjt_out  XM_bjt_out_0
timestamp 1662830870
transform 1 0 -1980 0 1 6780
box 0 0 6492 3916
use XM_feedbackmir2  XM_feedbackmir2_0
timestamp 1662719914
transform 1 0 -10768 0 1 9846
box -140 -160 2080 1600
use XM_feedbackmir  XM_feedbackmir_0
timestamp 1662675866
transform 1 0 -13500 0 1 8386
box -700 -500 2900 3100
use XM_otabias_nmos  XM_otabias_nmos_0
timestamp 1662818991
transform 1 0 -10166 0 1 7710
box -53 -53 1339 1105
use XM_otabias_pmos  XM_otabias_pmos_0
timestamp 1662818872
transform 1 0 -10817 0 1 8939
box -53 -53 1571 879
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662816987
transform 1 0 26563 0 1 -3003
box -17600 -7400 35500 15000
use XM_pdn  XM_pdn_0
timestamp 1662820526
transform 1 0 -8785 0 1 9133
box -53 -718 5502 1206
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662836520
transform 1 0 -8840 0 1 1874
box -5380 594 6776 6403
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_1
timestamp 1662836520
transform 1 0 -8840 0 1 -4044
box -5380 594 6776 6403
use sky130_fd_pr__res_high_po_1p41_6ZUZ5C  sky130_fd_pr__res_high_po_1p41_6ZUZ5C_0
timestamp 1662820359
transform 1 0 -8623 0 1 7103
box -307 -1408 307 1408
use sky130_fd_pr__res_high_po_1p41_GWJZ59  sky130_fd_pr__res_high_po_1p41_GWJZ59_0
timestamp 1662827202
transform 0 1 -3232 -1 0 -3669
box -307 -10998 307 10998
use sky130_fd_pr__res_high_po_1p41_HX7ZEK  sky130_fd_pr__res_high_po_1p41_HX7ZEK_0
timestamp 1662827686
transform 0 1 3187 -1 0 -3015
box -307 -5348 307 5348
use sky130_fd_pr__res_high_po_1p41_S8KB58  sky130_fd_pr__res_high_po_1p41_S8KB58_0
timestamp 1662758895
transform 0 1 -3253 -1 0 11177
box -307 -4837 307 4837
<< labels >>
flabel metal2 -9540 5700 -9480 7680 0 FreeSans 800 0 0 0 vb
flabel metal2 -11280 2300 1400 2500 0 FreeSans 1600 0 0 0 va
flabel metal3 -8760 8740 -8200 8840 0 FreeSans 800 0 0 0 vgate
<< end >>
