magic
tech sky130A
magscale 1 2
timestamp 1662323637
<< metal1 >>
rect 510 2600 520 2660
rect 580 2600 590 2660
rect 6290 1100 6300 1400
rect 6500 1100 6510 1400
rect 3346 966 3356 1031
rect 3338 928 3356 966
rect 3431 963 3441 1031
rect 3431 928 3459 963
rect 3338 907 3459 928
<< via1 >>
rect 520 2600 580 2660
rect 6300 1100 6500 1400
rect 3356 928 3431 1031
<< metal2 >>
rect 300 3670 650 3800
rect 280 2913 736 3045
rect -3780 2660 -3710 2670
rect -3780 2590 -3710 2600
rect -2480 2660 590 2670
rect -2480 2600 -1740 2660
rect -1670 2600 520 2660
rect 580 2600 590 2660
rect -2480 2590 590 2600
rect -4080 2330 -4000 2340
rect -4080 2260 -4000 2270
rect 301 2157 647 2289
rect 305 1401 651 1533
rect 6300 1400 6500 1410
rect 6300 1090 6500 1100
rect 3009 1031 3459 1047
rect 3009 928 3356 1031
rect 3431 928 3459 1031
rect 3009 907 3459 928
<< via2 >>
rect -3780 2600 -3710 2660
rect -1740 2600 -1670 2660
rect -4080 2270 -4000 2330
rect 6300 1100 6500 1400
<< metal3 >>
rect -1750 4874 -1740 4950
rect -1664 4874 -1654 4950
rect -3832 2665 -3702 4230
rect -3832 2660 -3700 2665
rect -3832 2600 -3780 2660
rect -3710 2600 -3700 2660
rect -3832 2595 -3700 2600
rect -1772 2660 -1642 4038
rect -1772 2600 -1740 2660
rect -1670 2600 -1642 2660
rect -3832 2590 -3702 2595
rect -1772 2560 -1642 2600
rect -4090 2330 -3990 2335
rect -4090 2270 -4080 2330
rect -4000 2270 -3990 2330
rect -4090 2265 -3990 2270
rect 6300 1405 6500 1800
rect 6290 1400 6510 1405
rect 6290 1100 6300 1400
rect 6500 1100 6510 1400
rect 6290 1095 6510 1100
<< via3 >>
rect -1740 4874 -1664 4950
<< metal4 >>
rect -1741 4950 -1663 4951
rect -1741 4874 -1740 4950
rect -1664 4940 -1663 4950
rect -1664 4880 3520 4940
rect -1664 4874 -1663 4880
rect -1741 4873 -1663 4874
use XM_actload2  XM_actload2_0
timestamp 1661870098
transform 1 0 -2047 0 1 753
box -53 -53 2571 3173
use XM_cs  XM_cs_0
timestamp 1662320303
transform 1 0 664 0 1 753
box -140 -53 2482 5609
use XM_diffpair  XM_diffpair_0
timestamp 1662313712
transform 1 0 -3688 0 1 2162
box -400 -1642 1600 1820
use XM_ppair  XM_ppair_0
timestamp 1662231221
transform 1 0 -5102 0 1 5030
box -220 -1160 4440 828
use XM_tail  XM_tail_0
timestamp 1662314158
transform 1 0 -5225 0 1 839
box -53 -51 1200 2931
use sky130_fd_pr__cap_mim_m3_1_EN3Q86  sky130_fd_pr__cap_mim_m3_1_EN3Q86_0
timestamp 1662322327
transform 1 0 4943 0 1 3949
box -1750 -2240 1647 2240
use sky130_fd_pr__res_high_po_2p85_7J2RPB  sky130_fd_pr__res_high_po_2p85_7J2RPB_0
timestamp 1662230297
transform 0 1 4968 -1 0 1241
box -451 -1808 451 1808
<< end >>
