magic
tech sky130A
magscale 1 2
timestamp 1662058138
<< metal1 >>
rect 750 370 760 460
rect 870 370 880 460
rect 1270 370 1280 460
rect 1390 370 1400 460
rect 2340 448 2386 460
rect 1316 360 1322 370
rect 1356 360 1362 370
rect 2340 150 2346 448
rect 2380 150 2386 448
rect 2598 448 2644 460
rect 240 60 250 150
rect 360 60 370 150
rect 1790 60 1800 150
rect 1910 60 1920 150
rect 2300 60 2310 150
rect 2420 60 2430 150
rect 2598 72 2604 448
rect 2638 72 2644 448
rect 2810 370 2820 460
rect 2930 370 2940 460
rect 3330 380 3340 470
rect 3450 380 3460 470
rect 3630 458 3676 470
rect 3372 370 3382 380
rect 3412 370 3422 380
rect 2598 60 2644 72
rect 2856 72 2862 370
rect 2896 72 2902 370
rect 2856 60 2902 72
rect 3372 82 3378 370
rect 3412 82 3418 370
rect 3372 70 3418 82
rect 3630 82 3636 458
rect 3670 82 3676 458
rect 3888 458 3934 470
rect 3888 160 3894 458
rect 3928 160 3934 458
rect 3630 70 3676 82
rect 3850 70 3860 160
rect 3970 70 3980 160
rect 70 -30 4140 20
rect 70 -360 4140 -310
rect 240 -480 250 -390
rect 360 -480 370 -390
rect 540 -402 586 -390
rect 282 -490 292 -480
rect 322 -490 332 -480
rect 282 -778 288 -490
rect 322 -778 328 -490
rect 282 -790 328 -778
rect 540 -778 546 -402
rect 580 -778 586 -402
rect 798 -402 844 -390
rect 798 -700 804 -402
rect 838 -700 844 -402
rect 1310 -412 1356 -400
rect 540 -790 586 -778
rect 760 -790 770 -700
rect 880 -790 890 -700
rect 1310 -710 1316 -412
rect 1350 -710 1356 -412
rect 1568 -412 1614 -400
rect 1270 -800 1280 -710
rect 1390 -800 1400 -710
rect 1568 -788 1574 -412
rect 1608 -788 1614 -412
rect 1780 -490 1790 -400
rect 1900 -490 1910 -400
rect 2300 -480 2310 -390
rect 2420 -480 2430 -390
rect 2600 -402 2646 -390
rect 2342 -490 2352 -480
rect 2382 -490 2392 -480
rect 1568 -800 1614 -788
rect 1826 -788 1832 -490
rect 1866 -788 1872 -490
rect 1826 -800 1872 -788
rect 2342 -778 2348 -490
rect 2382 -778 2388 -490
rect 2342 -790 2388 -778
rect 2600 -778 2606 -402
rect 2640 -778 2646 -402
rect 2858 -402 2904 -390
rect 2858 -700 2864 -402
rect 2898 -700 2904 -402
rect 3370 -422 3416 -410
rect 2600 -790 2646 -778
rect 2820 -790 2830 -700
rect 2940 -790 2950 -700
rect 3370 -720 3376 -422
rect 3410 -720 3416 -422
rect 3628 -422 3674 -410
rect 3330 -810 3340 -720
rect 3450 -810 3460 -720
rect 3628 -798 3634 -422
rect 3668 -798 3674 -422
rect 3840 -500 3850 -410
rect 3960 -500 3970 -410
rect 3628 -810 3674 -798
rect 3886 -798 3892 -500
rect 3926 -798 3932 -500
rect 3886 -810 3932 -798
<< via1 >>
rect 760 370 870 460
rect 1280 370 1390 460
rect 250 60 360 150
rect 1800 60 1910 150
rect 2310 60 2420 150
rect 2820 370 2930 460
rect 3340 380 3450 470
rect 3860 70 3970 160
rect 250 -480 360 -390
rect 770 -790 880 -700
rect 1280 -800 1390 -710
rect 1790 -490 1900 -400
rect 2310 -480 2420 -390
rect 2830 -790 2940 -700
rect 3340 -810 3450 -720
rect 3850 -500 3960 -410
<< metal2 >>
rect 750 470 3460 480
rect 750 460 3340 470
rect 750 370 760 460
rect 870 370 1280 460
rect 1390 370 2820 460
rect 2930 380 3340 460
rect 3450 380 3460 470
rect 2930 370 3460 380
rect 750 360 3460 370
rect 240 160 3980 170
rect 240 150 3860 160
rect 240 60 250 150
rect 360 60 1800 150
rect 1910 60 2310 150
rect 2420 70 3860 150
rect 3970 70 3980 160
rect 2420 60 3980 70
rect 240 50 3980 60
rect 250 -390 360 -380
rect 2310 -390 2420 -380
rect 240 -480 250 -390
rect 360 -400 2310 -390
rect 360 -480 1790 -400
rect 240 -490 1790 -480
rect 1900 -480 2310 -400
rect 2420 -410 3970 -390
rect 2420 -480 3850 -410
rect 1900 -490 3850 -480
rect 1790 -500 1900 -490
rect 3960 -490 3970 -410
rect 3850 -510 3960 -500
rect 770 -700 880 -690
rect 2830 -700 2940 -690
rect 760 -790 770 -710
rect 1280 -710 1390 -700
rect 880 -790 1280 -710
rect 760 -800 1280 -790
rect 1390 -790 2830 -710
rect 2940 -720 3460 -710
rect 2940 -790 3340 -720
rect 1390 -800 3340 -790
rect 760 -810 3340 -800
rect 3450 -810 3460 -720
rect 3340 -820 3450 -810
use sky130_fd_pr__pfet_01v8_lvt_B64SAM *sky130_fd_pr__pfet_01v8_lvt_B64SAM_0
timestamp 1661909013
transform 1 0 2109 0 1 224
box -2129 -264 2129 298
use sky130_fd_pr__pfet_01v8_lvt_MBDTEX  sky130_fd_pr__pfet_01v8_lvt_MBDTEX_0
timestamp 1661909182
transform 1 0 2109 0 1 -562
box -2129 -298 2129 264
<< labels >>
flabel space 220 -1160 380 -980 0 FreeSans 1600 0 0 0 B
flabel space 720 -1160 880 -980 0 FreeSans 1600 0 0 0 A
flabel space 1240 -1160 1400 -980 0 FreeSans 1600 0 0 0 A
flabel space 1760 -1160 1920 -980 0 FreeSans 1600 0 0 0 B
flabel space 2280 -1160 2440 -980 0 FreeSans 1600 0 0 0 B
flabel space 2780 -1160 2940 -980 0 FreeSans 1600 0 0 0 A
flabel space 3300 -1160 3460 -980 0 FreeSans 1600 0 0 0 A
flabel space 3820 -1160 3980 -980 0 FreeSans 1600 0 0 0 B
flabel space 240 648 400 828 0 FreeSans 1600 0 0 0 A
flabel space 740 648 900 828 0 FreeSans 1600 0 0 0 B
flabel space 1260 648 1420 828 0 FreeSans 1600 0 0 0 B
flabel space 1760 648 1920 828 0 FreeSans 1600 0 0 0 A
flabel space 2280 648 2440 828 0 FreeSans 1600 0 0 0 A
flabel space 2800 648 2960 828 0 FreeSans 1600 0 0 0 B
flabel space 3320 648 3480 828 0 FreeSans 1600 0 0 0 B
flabel space 3820 648 3980 828 0 FreeSans 1600 0 0 0 A
<< end >>
