magic
tech sky130A
magscale 1 2
timestamp 1662306324
<< locali >>
rect -20 2710 130 2790
rect 1010 2710 1160 2790
rect -20 2150 130 2230
rect 1010 2150 1160 2230
rect -20 1600 130 1680
rect 1010 1590 1160 1670
rect -20 1040 130 1120
rect 1010 1040 1160 1120
rect -20 480 130 560
rect 1010 480 1160 560
<< metal1 >>
rect 530 2550 540 2610
rect 610 2550 620 2610
rect 330 80 370 2350
rect 537 2305 607 2351
rect 530 2000 540 2060
rect 610 2000 620 2060
rect 537 1749 607 1795
rect 530 1430 540 1490
rect 610 1430 620 1490
rect 537 1193 607 1239
rect 530 870 540 930
rect 610 870 620 930
rect 537 637 607 683
rect 530 330 540 390
rect 610 330 620 390
rect 537 81 607 127
rect 780 80 820 2350
<< via1 >>
rect 540 2550 610 2610
rect 540 2000 610 2060
rect 540 1430 610 1490
rect 540 870 610 930
rect 540 330 610 390
<< metal2 >>
rect 540 2610 610 2620
rect 540 2060 610 2550
rect 540 1490 610 2000
rect 610 1430 1200 1490
rect 540 930 610 1430
rect 540 390 610 870
rect 540 320 610 330
use sky130_fd_pr__nfet_01v8_lvt_7MFZYU  sky130_fd_pr__nfet_01v8_lvt_7MFZYU_0
timestamp 1662302892
transform 1 0 572 0 1 1440
box -625 -1491 625 1491
<< end >>
