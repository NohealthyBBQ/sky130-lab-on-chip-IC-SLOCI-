magic
tech sky130A
magscale 1 2
timestamp 1662486269
<< pwell >>
rect -396 -7373 396 7373
<< nmoslvt >>
rect -200 5563 200 7163
rect -200 3745 200 5345
rect -200 1927 200 3527
rect -200 109 200 1709
rect -200 -1709 200 -109
rect -200 -3527 200 -1927
rect -200 -5345 200 -3745
rect -200 -7163 200 -5563
<< ndiff >>
rect -258 7151 -200 7163
rect -258 5575 -246 7151
rect -212 5575 -200 7151
rect -258 5563 -200 5575
rect 200 7151 258 7163
rect 200 5575 212 7151
rect 246 5575 258 7151
rect 200 5563 258 5575
rect -258 5333 -200 5345
rect -258 3757 -246 5333
rect -212 3757 -200 5333
rect -258 3745 -200 3757
rect 200 5333 258 5345
rect 200 3757 212 5333
rect 246 3757 258 5333
rect 200 3745 258 3757
rect -258 3515 -200 3527
rect -258 1939 -246 3515
rect -212 1939 -200 3515
rect -258 1927 -200 1939
rect 200 3515 258 3527
rect 200 1939 212 3515
rect 246 1939 258 3515
rect 200 1927 258 1939
rect -258 1697 -200 1709
rect -258 121 -246 1697
rect -212 121 -200 1697
rect -258 109 -200 121
rect 200 1697 258 1709
rect 200 121 212 1697
rect 246 121 258 1697
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -1697 -246 -121
rect -212 -1697 -200 -121
rect -258 -1709 -200 -1697
rect 200 -121 258 -109
rect 200 -1697 212 -121
rect 246 -1697 258 -121
rect 200 -1709 258 -1697
rect -258 -1939 -200 -1927
rect -258 -3515 -246 -1939
rect -212 -3515 -200 -1939
rect -258 -3527 -200 -3515
rect 200 -1939 258 -1927
rect 200 -3515 212 -1939
rect 246 -3515 258 -1939
rect 200 -3527 258 -3515
rect -258 -3757 -200 -3745
rect -258 -5333 -246 -3757
rect -212 -5333 -200 -3757
rect -258 -5345 -200 -5333
rect 200 -3757 258 -3745
rect 200 -5333 212 -3757
rect 246 -5333 258 -3757
rect 200 -5345 258 -5333
rect -258 -5575 -200 -5563
rect -258 -7151 -246 -5575
rect -212 -7151 -200 -5575
rect -258 -7163 -200 -7151
rect 200 -5575 258 -5563
rect 200 -7151 212 -5575
rect 246 -7151 258 -5575
rect 200 -7163 258 -7151
<< ndiffc >>
rect -246 5575 -212 7151
rect 212 5575 246 7151
rect -246 3757 -212 5333
rect 212 3757 246 5333
rect -246 1939 -212 3515
rect 212 1939 246 3515
rect -246 121 -212 1697
rect 212 121 246 1697
rect -246 -1697 -212 -121
rect 212 -1697 246 -121
rect -246 -3515 -212 -1939
rect 212 -3515 246 -1939
rect -246 -5333 -212 -3757
rect 212 -5333 246 -3757
rect -246 -7151 -212 -5575
rect 212 -7151 246 -5575
<< psubdiff >>
rect -360 7303 -264 7337
rect 264 7303 360 7337
rect -360 7241 -326 7303
rect 326 7241 360 7303
rect -360 -7303 -326 -7241
rect 326 -7303 360 -7241
rect -360 -7337 -264 -7303
rect 264 -7337 360 -7303
<< psubdiffcont >>
rect -264 7303 264 7337
rect -360 -7241 -326 7241
rect 326 -7241 360 7241
rect -264 -7337 264 -7303
<< poly >>
rect -200 7235 200 7251
rect -200 7201 -184 7235
rect 184 7201 200 7235
rect -200 7163 200 7201
rect -200 5525 200 5563
rect -200 5491 -184 5525
rect 184 5491 200 5525
rect -200 5475 200 5491
rect -200 5417 200 5433
rect -200 5383 -184 5417
rect 184 5383 200 5417
rect -200 5345 200 5383
rect -200 3707 200 3745
rect -200 3673 -184 3707
rect 184 3673 200 3707
rect -200 3657 200 3673
rect -200 3599 200 3615
rect -200 3565 -184 3599
rect 184 3565 200 3599
rect -200 3527 200 3565
rect -200 1889 200 1927
rect -200 1855 -184 1889
rect 184 1855 200 1889
rect -200 1839 200 1855
rect -200 1781 200 1797
rect -200 1747 -184 1781
rect 184 1747 200 1781
rect -200 1709 200 1747
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -1747 200 -1709
rect -200 -1781 -184 -1747
rect 184 -1781 200 -1747
rect -200 -1797 200 -1781
rect -200 -1855 200 -1839
rect -200 -1889 -184 -1855
rect 184 -1889 200 -1855
rect -200 -1927 200 -1889
rect -200 -3565 200 -3527
rect -200 -3599 -184 -3565
rect 184 -3599 200 -3565
rect -200 -3615 200 -3599
rect -200 -3673 200 -3657
rect -200 -3707 -184 -3673
rect 184 -3707 200 -3673
rect -200 -3745 200 -3707
rect -200 -5383 200 -5345
rect -200 -5417 -184 -5383
rect 184 -5417 200 -5383
rect -200 -5433 200 -5417
rect -200 -5491 200 -5475
rect -200 -5525 -184 -5491
rect 184 -5525 200 -5491
rect -200 -5563 200 -5525
rect -200 -7201 200 -7163
rect -200 -7235 -184 -7201
rect 184 -7235 200 -7201
rect -200 -7251 200 -7235
<< polycont >>
rect -184 7201 184 7235
rect -184 5491 184 5525
rect -184 5383 184 5417
rect -184 3673 184 3707
rect -184 3565 184 3599
rect -184 1855 184 1889
rect -184 1747 184 1781
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -1781 184 -1747
rect -184 -1889 184 -1855
rect -184 -3599 184 -3565
rect -184 -3707 184 -3673
rect -184 -5417 184 -5383
rect -184 -5525 184 -5491
rect -184 -7235 184 -7201
<< locali >>
rect -360 7303 -264 7337
rect 264 7303 360 7337
rect -360 7241 -326 7303
rect 326 7241 360 7303
rect -200 7201 -184 7235
rect 184 7201 200 7235
rect -246 7151 -212 7167
rect -246 5559 -212 5575
rect 212 7151 246 7167
rect 212 5559 246 5575
rect -200 5491 -184 5525
rect 184 5491 200 5525
rect -200 5383 -184 5417
rect 184 5383 200 5417
rect -246 5333 -212 5349
rect -246 3741 -212 3757
rect 212 5333 246 5349
rect 212 3741 246 3757
rect -200 3673 -184 3707
rect 184 3673 200 3707
rect -200 3565 -184 3599
rect 184 3565 200 3599
rect -246 3515 -212 3531
rect -246 1923 -212 1939
rect 212 3515 246 3531
rect 212 1923 246 1939
rect -200 1855 -184 1889
rect 184 1855 200 1889
rect -200 1747 -184 1781
rect 184 1747 200 1781
rect -246 1697 -212 1713
rect -246 105 -212 121
rect 212 1697 246 1713
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -1713 -212 -1697
rect 212 -121 246 -105
rect 212 -1713 246 -1697
rect -200 -1781 -184 -1747
rect 184 -1781 200 -1747
rect -200 -1889 -184 -1855
rect 184 -1889 200 -1855
rect -246 -1939 -212 -1923
rect -246 -3531 -212 -3515
rect 212 -1939 246 -1923
rect 212 -3531 246 -3515
rect -200 -3599 -184 -3565
rect 184 -3599 200 -3565
rect -200 -3707 -184 -3673
rect 184 -3707 200 -3673
rect -246 -3757 -212 -3741
rect -246 -5349 -212 -5333
rect 212 -3757 246 -3741
rect 212 -5349 246 -5333
rect -200 -5417 -184 -5383
rect 184 -5417 200 -5383
rect -200 -5525 -184 -5491
rect 184 -5525 200 -5491
rect -246 -5575 -212 -5559
rect -246 -7167 -212 -7151
rect 212 -5575 246 -5559
rect 212 -7167 246 -7151
rect -200 -7235 -184 -7201
rect 184 -7235 200 -7201
rect -360 -7303 -326 -7241
rect 326 -7303 360 -7241
rect -360 -7337 -264 -7303
rect 264 -7337 360 -7303
<< viali >>
rect -184 7201 184 7235
rect -246 5575 -212 7151
rect 212 5575 246 7151
rect -184 5491 184 5525
rect -184 5383 184 5417
rect -246 3757 -212 5333
rect 212 3757 246 5333
rect -184 3673 184 3707
rect -184 3565 184 3599
rect -246 1939 -212 3515
rect 212 1939 246 3515
rect -184 1855 184 1889
rect -184 1747 184 1781
rect -246 121 -212 1697
rect 212 121 246 1697
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -1697 -212 -121
rect 212 -1697 246 -121
rect -184 -1781 184 -1747
rect -184 -1889 184 -1855
rect -246 -3515 -212 -1939
rect 212 -3515 246 -1939
rect -184 -3599 184 -3565
rect -184 -3707 184 -3673
rect -246 -5333 -212 -3757
rect 212 -5333 246 -3757
rect -184 -5417 184 -5383
rect -184 -5525 184 -5491
rect -246 -7151 -212 -5575
rect 212 -7151 246 -5575
rect -184 -7235 184 -7201
<< metal1 >>
rect -196 7235 196 7241
rect -196 7201 -184 7235
rect 184 7201 196 7235
rect -196 7195 196 7201
rect -252 7151 -206 7163
rect -252 5575 -246 7151
rect -212 5575 -206 7151
rect -252 5563 -206 5575
rect 206 7151 252 7163
rect 206 5575 212 7151
rect 246 5575 252 7151
rect 206 5563 252 5575
rect -196 5525 196 5531
rect -196 5491 -184 5525
rect 184 5491 196 5525
rect -196 5485 196 5491
rect -196 5417 196 5423
rect -196 5383 -184 5417
rect 184 5383 196 5417
rect -196 5377 196 5383
rect -252 5333 -206 5345
rect -252 3757 -246 5333
rect -212 3757 -206 5333
rect -252 3745 -206 3757
rect 206 5333 252 5345
rect 206 3757 212 5333
rect 246 3757 252 5333
rect 206 3745 252 3757
rect -196 3707 196 3713
rect -196 3673 -184 3707
rect 184 3673 196 3707
rect -196 3667 196 3673
rect -196 3599 196 3605
rect -196 3565 -184 3599
rect 184 3565 196 3599
rect -196 3559 196 3565
rect -252 3515 -206 3527
rect -252 1939 -246 3515
rect -212 1939 -206 3515
rect -252 1927 -206 1939
rect 206 3515 252 3527
rect 206 1939 212 3515
rect 246 1939 252 3515
rect 206 1927 252 1939
rect -196 1889 196 1895
rect -196 1855 -184 1889
rect 184 1855 196 1889
rect -196 1849 196 1855
rect -196 1781 196 1787
rect -196 1747 -184 1781
rect 184 1747 196 1781
rect -196 1741 196 1747
rect -252 1697 -206 1709
rect -252 121 -246 1697
rect -212 121 -206 1697
rect -252 109 -206 121
rect 206 1697 252 1709
rect 206 121 212 1697
rect 246 121 252 1697
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -1697 -246 -121
rect -212 -1697 -206 -121
rect -252 -1709 -206 -1697
rect 206 -121 252 -109
rect 206 -1697 212 -121
rect 246 -1697 252 -121
rect 206 -1709 252 -1697
rect -196 -1747 196 -1741
rect -196 -1781 -184 -1747
rect 184 -1781 196 -1747
rect -196 -1787 196 -1781
rect -196 -1855 196 -1849
rect -196 -1889 -184 -1855
rect 184 -1889 196 -1855
rect -196 -1895 196 -1889
rect -252 -1939 -206 -1927
rect -252 -3515 -246 -1939
rect -212 -3515 -206 -1939
rect -252 -3527 -206 -3515
rect 206 -1939 252 -1927
rect 206 -3515 212 -1939
rect 246 -3515 252 -1939
rect 206 -3527 252 -3515
rect -196 -3565 196 -3559
rect -196 -3599 -184 -3565
rect 184 -3599 196 -3565
rect -196 -3605 196 -3599
rect -196 -3673 196 -3667
rect -196 -3707 -184 -3673
rect 184 -3707 196 -3673
rect -196 -3713 196 -3707
rect -252 -3757 -206 -3745
rect -252 -5333 -246 -3757
rect -212 -5333 -206 -3757
rect -252 -5345 -206 -5333
rect 206 -3757 252 -3745
rect 206 -5333 212 -3757
rect 246 -5333 252 -3757
rect 206 -5345 252 -5333
rect -196 -5383 196 -5377
rect -196 -5417 -184 -5383
rect 184 -5417 196 -5383
rect -196 -5423 196 -5417
rect -196 -5491 196 -5485
rect -196 -5525 -184 -5491
rect 184 -5525 196 -5491
rect -196 -5531 196 -5525
rect -252 -5575 -206 -5563
rect -252 -7151 -246 -5575
rect -212 -7151 -206 -5575
rect -252 -7163 -206 -7151
rect 206 -5575 252 -5563
rect 206 -7151 212 -5575
rect 246 -7151 252 -5575
rect 206 -7163 252 -7151
rect -196 -7201 196 -7195
rect -196 -7235 -184 -7201
rect 184 -7235 196 -7201
rect -196 -7241 196 -7235
<< properties >>
string FIXED_BBOX -343 -7320 343 7320
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8.0 l 2.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
