magic
tech sky130A
magscale 1 2
timestamp 1662978535
<< metal1 >>
rect 1220 8010 1230 8074
rect 1294 8010 1304 8074
rect 230 3470 270 6820
rect 4880 5730 20600 5770
rect 230 3430 1500 3470
rect 1460 3040 1500 3430
rect 4750 3410 4780 4510
rect 3450 3380 4780 3410
rect 3450 2820 3480 3380
rect 3450 2790 3570 2820
rect 20560 2300 20600 5730
rect 110 1770 4650 1800
rect 110 1710 4150 1740
rect 4120 1510 4150 1710
rect 19936 1700 23570 1738
rect 19936 1592 19978 1700
rect 17752 1558 19978 1592
rect 5550 1510 5580 1520
rect 4120 1480 5580 1510
rect 3510 628 3570 658
rect 1460 60 1500 422
rect 280 20 1500 60
rect 280 -2310 320 20
rect 1250 -810 1260 -700
rect 1370 -810 1380 -700
rect 3510 -3630 3540 628
rect 21490 -1740 21520 1180
rect 4930 -1770 21520 -1740
rect 3510 -3660 4870 -3630
rect 4840 -4250 4870 -3660
<< via1 >>
rect 1230 8010 1294 8074
rect 1260 -810 1370 -700
<< metal2 >>
rect 1230 8074 1294 8084
rect 1230 8000 1294 8010
rect 710 4314 774 4324
rect 710 4240 774 4250
rect 2256 3416 2376 4718
rect 720 -556 784 -546
rect 720 -630 784 -620
rect 730 -1030 770 -630
rect 1260 -700 1370 -690
rect 2300 -810 2420 10
rect 1260 -820 1370 -810
<< via2 >>
rect 1230 8010 1294 8074
rect 710 4250 774 4314
rect 720 -620 784 -556
rect 1260 -810 1370 -700
<< metal3 >>
rect 1220 8074 1330 8110
rect 1220 8010 1230 8074
rect 1294 8010 1330 8074
rect 1220 8000 1330 8010
rect 690 4314 800 4330
rect 286 2994 426 4259
rect 690 4250 710 4314
rect 774 4250 800 4314
rect 690 4240 800 4250
rect 330 -812 470 453
rect 710 -556 800 -530
rect 710 -620 720 -556
rect 784 -620 800 -556
rect 710 -660 800 -620
rect 1250 -700 1380 -695
rect 1250 -810 1260 -700
rect 1370 -810 1380 -700
rect 1250 -815 1380 -810
<< via3 >>
rect 1230 8010 1294 8074
rect 710 4250 774 4314
rect 720 -620 784 -556
rect 1260 -810 1370 -700
<< metal4 >>
rect 1260 8075 1330 8110
rect 1229 8074 1330 8075
rect 1229 8010 1230 8074
rect 1294 8010 1330 8074
rect 1229 8009 1330 8010
rect 709 4314 775 4315
rect 709 4250 710 4314
rect 774 4260 775 4314
rect 774 4250 790 4260
rect 709 4249 790 4250
rect 710 -556 790 4249
rect 710 -620 720 -556
rect 784 -620 790 -556
rect 710 -630 790 -620
rect 1260 -699 1330 8009
rect 1259 -700 1371 -699
rect 1259 -810 1260 -700
rect 1370 -810 1371 -700
rect 1259 -811 1371 -810
use cmfb1  cmfb1_0
timestamp 1662938211
transform 0 1 8026 -1 0 697
box -8100 -7760 -2801 18240
use cmfb1  cmfb1_1
timestamp 1662938211
transform 0 1 8070 -1 0 -8125
box -8100 -7760 -2801 18240
use cons_cw  cons_cw_0
timestamp 1662976792
transform 1 0 -46324 0 1 8198
box 46324 -8198 69992 -4736
<< labels >>
rlabel space 416 0 23486 390 0 vdd
rlabel space 330 -1255 470 688 0 vss
rlabel metal1 230 3430 270 6820 0 vout2p
rlabel metal1 20560 2890 20600 5770 0 vout2n
rlabel metal1 280 -2310 320 60 0 vd21
rlabel metal1 21490 -1770 21520 570 0 vd22
rlabel space 686 7777 726 8207 0 vbias2
rlabel metal1 3450 2790 3480 3410 0 vo22
rlabel metal1 3510 -3660 3540 658 0 vo21
rlabel metal1 110 1710 4150 1740 0 vout1p
rlabel metal3 1220 8074 1330 8110 0 vref
rlabel space 110 1770 4696 1800 0 vc
rlabel metal1 19936 1700 23570 1738 0 vout1n
<< end >>
