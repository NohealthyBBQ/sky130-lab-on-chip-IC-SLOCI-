magic
tech sky130A
magscale 1 2
timestamp 1662769262
<< metal1 >>
rect -10 860 0 920
rect 60 860 70 920
rect 450 860 460 920
rect 520 860 530 920
rect 910 860 920 920
rect 980 860 990 920
rect 1370 860 1380 920
rect 1440 860 1450 920
rect 1830 860 1840 920
rect 1900 860 1910 920
rect 62 -98 1828 56
rect -10 -960 0 -900
rect 60 -960 70 -900
rect 450 -960 460 -900
rect 520 -960 530 -900
rect 910 -960 920 -900
rect 980 -960 990 -900
rect 1370 -960 1380 -900
rect 1440 -960 1450 -900
rect 1830 -960 1840 -900
rect 1900 -960 1910 -900
rect -10 -2640 0 -2580
rect 60 -2640 70 -2580
rect 450 -2640 460 -2580
rect 520 -2640 530 -2580
rect 910 -2640 920 -2580
rect 980 -2640 990 -2580
rect 1370 -2640 1380 -2580
rect 1440 -2640 1450 -2580
rect 1830 -2640 1840 -2580
rect 1900 -2640 1910 -2580
rect 62 -3610 1828 -3456
rect -10 -4460 0 -4400
rect 60 -4460 70 -4400
rect 450 -4460 460 -4400
rect 520 -4460 530 -4400
rect 910 -4460 920 -4400
rect 980 -4460 990 -4400
rect 1370 -4460 1380 -4400
rect 1440 -4460 1450 -4400
rect 1830 -4460 1840 -4400
rect 1900 -4460 1910 -4400
<< via1 >>
rect 0 860 60 920
rect 460 860 520 920
rect 920 860 980 920
rect 1380 860 1440 920
rect 1840 860 1900 920
rect 0 -960 60 -900
rect 460 -960 520 -900
rect 920 -960 980 -900
rect 1380 -960 1440 -900
rect 1840 -960 1900 -900
rect 0 -2640 60 -2580
rect 460 -2640 520 -2580
rect 920 -2640 980 -2580
rect 1380 -2640 1440 -2580
rect 1840 -2640 1900 -2580
rect 0 -4460 60 -4400
rect 460 -4460 520 -4400
rect 920 -4460 980 -4400
rect 1380 -4460 1440 -4400
rect 1840 -4460 1900 -4400
<< metal2 >>
rect 0 1640 1900 1700
rect 0 920 60 1640
rect 0 -900 60 860
rect 0 -970 60 -960
rect 460 920 520 930
rect 460 -900 520 860
rect 460 -1746 520 -960
rect 920 920 980 1640
rect 920 -900 980 860
rect 920 -970 980 -960
rect 1380 920 1440 930
rect 1380 -900 1440 860
rect 1380 -1746 1440 -960
rect 1840 920 1900 1640
rect 1840 -900 1900 860
rect 1840 -970 1900 -960
rect 460 -1806 1440 -1746
rect 0 -2580 60 -2570
rect 0 -4400 60 -2640
rect 0 -5180 60 -4460
rect 460 -2580 520 -1806
rect 460 -4400 520 -2640
rect 460 -4470 520 -4460
rect 920 -2580 980 -2570
rect 920 -4400 980 -2640
rect 920 -5180 980 -4460
rect 1380 -2580 1440 -1806
rect 1380 -4400 1440 -2640
rect 1380 -4470 1440 -4460
rect 1840 -2580 1900 -2570
rect 1840 -4400 1900 -2640
rect 1840 -5180 1900 -4460
rect 0 -5240 1900 -5180
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_0
timestamp 1662766393
transform 1 0 945 0 1 -899
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_1
timestamp 1662766393
transform 1 0 945 0 1 -4411
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_0
timestamp 1662766393
transform 1 0 945 0 1 857
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_1
timestamp 1662766393
transform 1 0 945 0 1 -2655
box -945 -857 945 857
<< end >>
