magic
tech sky130A
magscale 1 2
timestamp 1662721300
<< metal1 >>
rect 70 680 80 740
rect 140 680 150 740
rect 590 680 600 740
rect 660 680 670 740
rect 1110 680 1120 740
rect 1180 680 1190 740
rect 330 520 340 580
rect 400 520 410 580
rect 850 520 860 580
rect 920 520 930 580
rect 1370 520 1380 580
rect 1440 520 1450 580
rect 144 448 1380 480
rect 70 320 80 380
rect 140 320 150 380
rect 590 320 600 380
rect 660 320 670 380
rect 330 160 340 220
rect 400 160 410 220
rect 740 119 780 448
rect 1110 320 1120 380
rect 1180 320 1190 380
rect 850 160 860 220
rect 920 160 930 220
rect 1370 160 1380 220
rect 1440 160 1450 220
rect 143 85 1367 119
rect 740 80 780 85
<< via1 >>
rect 80 680 140 740
rect 600 680 660 740
rect 1120 680 1180 740
rect 340 520 400 580
rect 860 520 920 580
rect 1380 520 1440 580
rect 80 320 140 380
rect 600 320 660 380
rect 340 160 400 220
rect 1120 320 1180 380
rect 860 160 920 220
rect 1380 160 1440 220
<< metal2 >>
rect 80 740 140 750
rect 600 740 660 750
rect 1120 740 1180 750
rect 140 680 600 740
rect 660 680 1120 740
rect 80 380 140 680
rect 600 670 660 680
rect 1120 670 1180 680
rect 340 580 400 590
rect 1380 580 1440 590
rect 400 520 860 580
rect 920 520 1380 580
rect 340 510 400 520
rect 600 380 660 390
rect 1120 380 1180 390
rect 140 320 600 380
rect 660 320 1120 380
rect 80 310 140 320
rect 600 310 660 320
rect 1120 310 1180 320
rect 340 220 400 230
rect 1380 220 1440 520
rect 400 160 860 220
rect 920 160 1380 220
rect 340 150 400 160
rect 1380 150 1440 160
use sky130_fd_pr__pfet_01v8_lvt_9UVN44  sky130_fd_pr__pfet_01v8_lvt_9UVN44_0
timestamp 1662720466
transform 1 0 759 0 1 413
box -812 -466 812 466
<< end >>
