** sch_path: /foss/designs/sumprj/hiarachy_final/cap_bank.sch
.subckt cap_bank IN GND ctrll1 ctrll2 ctrll3 ctrll4 ctrll5
*.PININFO IN:I GND:I ctrll1:I ctrll2:I ctrll3:I ctrll4:I ctrll5:I
XC6 IN net1 sky130_fd_pr__cap_mim_m3_2 W=2 L=2 VM=1 m=1
XC1 IN net5 sky130_fd_pr__cap_mim_m3_2 W=2 L=2 VM=1 m=1
XC2 IN net4 sky130_fd_pr__cap_mim_m3_2 W=3 L=2 VM=1 m=1
XC3 IN net3 sky130_fd_pr__cap_mim_m3_2 W=3 L=4 VM=1 m=1
XC4 IN net2 sky130_fd_pr__cap_mim_m3_2 W=6 L=4 VM=1 m=1
XM1 net1 ctrll1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net5 ctrll2 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net4 ctrll3 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 ctrll4 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 ctrll5 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends
.end
