magic
tech sky130A
magscale 1 2
timestamp 1662486269
<< pwell >>
rect -296 -2337 296 2337
<< nmoslvt >>
rect -100 1227 100 2127
rect -100 109 100 1009
rect -100 -1009 100 -109
rect -100 -2127 100 -1227
<< ndiff >>
rect -158 2115 -100 2127
rect -158 1239 -146 2115
rect -112 1239 -100 2115
rect -158 1227 -100 1239
rect 100 2115 158 2127
rect 100 1239 112 2115
rect 146 1239 158 2115
rect 100 1227 158 1239
rect -158 997 -100 1009
rect -158 121 -146 997
rect -112 121 -100 997
rect -158 109 -100 121
rect 100 997 158 1009
rect 100 121 112 997
rect 146 121 158 997
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -997 -146 -121
rect -112 -997 -100 -121
rect -158 -1009 -100 -997
rect 100 -121 158 -109
rect 100 -997 112 -121
rect 146 -997 158 -121
rect 100 -1009 158 -997
rect -158 -1239 -100 -1227
rect -158 -2115 -146 -1239
rect -112 -2115 -100 -1239
rect -158 -2127 -100 -2115
rect 100 -1239 158 -1227
rect 100 -2115 112 -1239
rect 146 -2115 158 -1239
rect 100 -2127 158 -2115
<< ndiffc >>
rect -146 1239 -112 2115
rect 112 1239 146 2115
rect -146 121 -112 997
rect 112 121 146 997
rect -146 -997 -112 -121
rect 112 -997 146 -121
rect -146 -2115 -112 -1239
rect 112 -2115 146 -1239
<< psubdiff >>
rect -260 2267 -164 2301
rect 164 2267 260 2301
rect -260 2205 -226 2267
rect 226 2205 260 2267
rect -260 -2267 -226 -2205
rect 226 -2267 260 -2205
rect -260 -2301 -164 -2267
rect 164 -2301 260 -2267
<< psubdiffcont >>
rect -164 2267 164 2301
rect -260 -2205 -226 2205
rect 226 -2205 260 2205
rect -164 -2301 164 -2267
<< poly >>
rect -100 2199 100 2215
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -100 2127 100 2165
rect -100 1189 100 1227
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1139 100 1155
rect -100 1081 100 1097
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -100 1009 100 1047
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1047 100 -1009
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1097 100 -1081
rect -100 -1155 100 -1139
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -100 -1227 100 -1189
rect -100 -2165 100 -2127
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2215 100 -2199
<< polycont >>
rect -84 2165 84 2199
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -84 -2199 84 -2165
<< locali >>
rect -260 2267 -164 2301
rect 164 2267 260 2301
rect -260 2205 -226 2267
rect 226 2205 260 2267
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -146 2115 -112 2131
rect -146 1223 -112 1239
rect 112 2115 146 2131
rect 112 1223 146 1239
rect -100 1155 -84 1189
rect 84 1155 100 1189
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -146 997 -112 1013
rect -146 105 -112 121
rect 112 997 146 1013
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1013 -112 -997
rect 112 -121 146 -105
rect 112 -1013 146 -997
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1189 -84 -1155
rect 84 -1189 100 -1155
rect -146 -1239 -112 -1223
rect -146 -2131 -112 -2115
rect 112 -1239 146 -1223
rect 112 -2131 146 -2115
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -260 -2267 -226 -2205
rect 226 -2267 260 -2205
rect -260 -2301 -164 -2267
rect 164 -2301 260 -2267
<< viali >>
rect -84 2165 84 2199
rect -146 1239 -112 2115
rect 112 1239 146 2115
rect -84 1155 84 1189
rect -84 1047 84 1081
rect -146 121 -112 997
rect 112 121 146 997
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -997 -112 -121
rect 112 -997 146 -121
rect -84 -1081 84 -1047
rect -84 -1189 84 -1155
rect -146 -2115 -112 -1239
rect 112 -2115 146 -1239
rect -84 -2199 84 -2165
<< metal1 >>
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect -152 2115 -106 2127
rect -152 1239 -146 2115
rect -112 1239 -106 2115
rect -152 1227 -106 1239
rect 106 2115 152 2127
rect 106 1239 112 2115
rect 146 1239 152 2115
rect 106 1227 152 1239
rect -96 1189 96 1195
rect -96 1155 -84 1189
rect 84 1155 96 1189
rect -96 1149 96 1155
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect -152 997 -106 1009
rect -152 121 -146 997
rect -112 121 -106 997
rect -152 109 -106 121
rect 106 997 152 1009
rect 106 121 112 997
rect 146 121 152 997
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -997 -146 -121
rect -112 -997 -106 -121
rect -152 -1009 -106 -997
rect 106 -121 152 -109
rect 106 -997 112 -121
rect 146 -997 152 -121
rect 106 -1009 152 -997
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
rect -96 -1155 96 -1149
rect -96 -1189 -84 -1155
rect 84 -1189 96 -1155
rect -96 -1195 96 -1189
rect -152 -1239 -106 -1227
rect -152 -2115 -146 -1239
rect -112 -2115 -106 -1239
rect -152 -2127 -106 -2115
rect 106 -1239 152 -1227
rect 106 -2115 112 -1239
rect 146 -2115 152 -1239
rect 106 -2127 152 -2115
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
<< properties >>
string FIXED_BBOX -243 -2284 243 2284
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.5 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
