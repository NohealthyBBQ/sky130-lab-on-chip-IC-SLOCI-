magic
tech sky130A
magscale 1 2
timestamp 1662494177
<< nwell >>
rect -4 1996 2272 3500
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_0
timestamp 1662493693
transform 1 0 284 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_1
timestamp 1662493693
transform 1 0 542 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_2
timestamp 1662493693
transform 1 0 800 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_3
timestamp 1662493693
transform 1 0 1058 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_4
timestamp 1662493693
transform 1 0 1316 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_5
timestamp 1662493693
transform 1 0 1574 0 1 2740
box -194 -712 194 745
use sky130_fd_pr__pfet_01v8_lvt_9UV3G5  sky130_fd_pr__pfet_01v8_lvt_9UV3G5_6
timestamp 1662493693
transform 1 0 1832 0 1 2740
box -194 -712 194 745
<< end >>
