magic
tech sky130A
magscale 1 2
timestamp 1662067076
<< nwell >>
rect -220 -1060 4440 720
<< nsubdiff >>
rect -140 580 520 640
rect 860 580 1300 640
rect 1640 580 2580 640
rect 2920 580 3360 640
rect 3700 580 4360 640
rect -140 460 -80 580
rect -140 -140 -80 60
rect 4300 460 4360 580
rect 4300 -140 4360 60
rect -140 -200 520 -140
rect 860 -200 1300 -140
rect 1640 -200 2580 -140
rect 2920 -200 3360 -140
rect 3700 -200 4360 -140
rect -140 -400 -80 -200
rect -140 -920 -80 -800
rect 4300 -400 4360 -200
rect 4300 -920 4360 -800
rect -140 -980 520 -920
rect 860 -980 1300 -920
rect 1640 -980 2580 -920
rect 2920 -980 3360 -920
rect 3700 -980 4360 -920
<< nsubdiffcont >>
rect 520 580 860 640
rect 1300 580 1640 640
rect 2580 580 2920 640
rect 3360 580 3700 640
rect -140 60 -80 460
rect 4300 60 4360 460
rect 520 -200 860 -140
rect 1300 -200 1640 -140
rect 2580 -200 2920 -140
rect 3360 -200 3700 -140
rect -140 -800 -80 -400
rect 4300 -800 4360 -400
rect 520 -980 860 -920
rect 1300 -980 1640 -920
rect 2580 -980 2920 -920
rect 3360 -980 3700 -920
<< locali >>
rect -140 580 520 640
rect 860 580 1300 640
rect 1640 580 2580 640
rect 2920 580 3360 640
rect 3700 580 4360 640
rect -140 460 -80 580
rect -140 -140 -80 60
rect 4300 460 4360 580
rect 4300 -140 4360 60
rect -140 -200 520 -140
rect 860 -200 1300 -140
rect 1640 -200 2580 -140
rect 2920 -200 3360 -140
rect 3700 -200 4360 -140
rect -140 -400 -80 -200
rect -140 -920 -80 -800
rect 4300 -400 4360 -200
rect 4300 -920 4360 -800
rect -140 -980 520 -920
rect 860 -980 1300 -920
rect 1640 -980 2580 -920
rect 2920 -980 3360 -920
rect 3700 -980 4360 -920
<< viali >>
rect 520 580 860 640
rect 1300 580 1640 640
rect 2580 580 2920 640
rect 3360 580 3700 640
rect 520 -980 860 -920
rect 1300 -980 1640 -920
rect 2580 -980 2920 -920
rect 3360 -980 3700 -920
<< metal1 >>
rect -140 640 4360 646
rect -140 580 520 640
rect 860 580 1300 640
rect 1640 580 2580 640
rect 2920 580 3360 640
rect 3700 580 4360 640
rect -140 574 4360 580
rect -140 -914 -80 574
rect 22 420 68 574
rect 538 420 584 574
rect 750 370 760 460
rect 870 370 880 460
rect 1054 420 1100 574
rect 1270 370 1280 460
rect 1390 370 1400 460
rect 1570 420 1616 574
rect 2086 420 2132 574
rect 2340 448 2386 460
rect 1316 360 1322 370
rect 1356 360 1362 370
rect 2340 150 2346 448
rect 2380 150 2386 448
rect 2598 448 2648 574
rect 240 60 250 150
rect 360 60 370 150
rect 1790 60 1800 150
rect 1910 60 1920 150
rect 2300 60 2310 150
rect 2420 60 2430 150
rect 2598 72 2604 448
rect 2810 370 2820 460
rect 2930 370 2940 460
rect 3118 449 3164 574
rect 3330 380 3340 470
rect 3450 380 3460 470
rect 3630 454 3680 574
rect 3888 459 3938 460
rect 3888 458 3934 459
rect 3372 370 3382 380
rect 3412 370 3422 380
rect 2856 72 2862 370
rect 2896 72 2902 370
rect 2598 60 2638 72
rect 2856 60 2902 72
rect 3372 82 3378 370
rect 3412 82 3418 370
rect 3372 70 3418 82
rect 3630 82 3636 454
rect 3670 82 3676 454
rect 3888 160 3894 458
rect 3928 160 3934 458
rect 4150 457 4196 574
rect 3630 70 3676 82
rect 3850 70 3860 160
rect 3970 70 3980 160
rect 280 20 330 60
rect 1830 20 1880 60
rect 2340 20 2390 60
rect 3890 20 3940 70
rect 70 -30 4140 20
rect 280 -310 330 -30
rect 1830 -310 1880 -30
rect 2340 -310 2390 -30
rect 3890 -310 3940 -30
rect 70 -360 4140 -310
rect 240 -480 250 -390
rect 360 -480 370 -390
rect 540 -402 586 -390
rect 282 -490 292 -480
rect 322 -490 332 -480
rect 282 -778 288 -490
rect 322 -778 328 -490
rect 21 -914 68 -789
rect 282 -790 328 -778
rect 540 -778 546 -402
rect 580 -778 586 -402
rect 798 -402 844 -390
rect 798 -700 804 -402
rect 838 -700 844 -402
rect 1310 -412 1356 -400
rect 540 -787 586 -778
rect 538 -914 586 -787
rect 760 -790 770 -700
rect 880 -790 890 -700
rect 1310 -710 1316 -412
rect 1350 -710 1356 -412
rect 1568 -412 1614 -400
rect 1054 -914 1100 -789
rect 1270 -800 1280 -710
rect 1390 -800 1400 -710
rect 1568 -788 1574 -412
rect 1608 -788 1614 -412
rect 1780 -490 1790 -400
rect 1900 -490 1910 -400
rect 2300 -480 2310 -390
rect 2420 -480 2430 -390
rect 2600 -402 2646 -390
rect 2342 -490 2352 -480
rect 2382 -490 2392 -480
rect 1568 -794 1614 -788
rect 1826 -788 1832 -490
rect 1866 -788 1872 -490
rect 1568 -914 1616 -794
rect 1826 -800 1872 -788
rect 2342 -778 2348 -490
rect 2382 -778 2388 -490
rect 2342 -790 2388 -778
rect 2600 -778 2606 -402
rect 2640 -778 2646 -402
rect 2858 -402 2904 -390
rect 2858 -700 2864 -402
rect 2898 -700 2904 -402
rect 3370 -422 3416 -410
rect 2600 -784 2646 -778
rect 2086 -914 2132 -794
rect 2600 -914 2648 -784
rect 2820 -790 2830 -700
rect 2940 -790 2950 -700
rect 3370 -720 3376 -422
rect 3410 -720 3416 -422
rect 3628 -422 3674 -410
rect 3118 -914 3164 -778
rect 3330 -810 3340 -720
rect 3450 -810 3460 -720
rect 3628 -782 3634 -422
rect 3668 -782 3674 -422
rect 3840 -500 3850 -410
rect 3960 -500 3970 -410
rect 3628 -914 3680 -782
rect 3886 -798 3892 -500
rect 3926 -798 3932 -500
rect 3886 -810 3932 -798
rect 4150 -914 4196 -775
rect 4300 -914 4360 574
rect -140 -920 4360 -914
rect -140 -980 520 -920
rect 860 -980 1300 -920
rect 1640 -980 2580 -920
rect 2920 -980 3360 -920
rect 3700 -980 4360 -920
rect -140 -986 4360 -980
<< via1 >>
rect 760 370 870 460
rect 1280 370 1390 460
rect 250 60 360 150
rect 1800 60 1910 150
rect 2310 60 2420 150
rect 2820 370 2930 460
rect 3340 380 3450 470
rect 3860 70 3970 160
rect 250 -480 360 -390
rect 770 -790 880 -700
rect 1280 -800 1390 -710
rect 1790 -490 1900 -400
rect 2310 -480 2420 -390
rect 2830 -790 2940 -700
rect 3340 -810 3450 -720
rect 3850 -500 3960 -410
<< metal2 >>
rect 750 470 3460 480
rect 750 460 3340 470
rect 3450 460 3460 470
rect 750 370 758 460
rect 870 370 1280 460
rect 1390 370 2820 460
rect 2930 370 3340 460
rect 3452 370 3460 460
rect 750 360 3460 370
rect 240 160 3980 170
rect 240 150 3860 160
rect 240 60 250 150
rect 360 60 1280 150
rect 1392 60 1800 150
rect 1910 60 2310 150
rect 2420 60 2830 150
rect 2942 70 3860 150
rect 3970 70 3980 160
rect 2942 60 3980 70
rect 240 50 3980 60
rect 250 -390 360 -380
rect 760 -390 872 -380
rect 2310 -390 2420 -380
rect 3340 -390 3452 -380
rect 240 -480 250 -390
rect 360 -480 760 -390
rect 872 -400 2310 -390
rect 872 -480 1790 -400
rect 240 -490 1790 -480
rect 1900 -480 2310 -400
rect 2420 -480 3340 -390
rect 3452 -410 3970 -390
rect 3452 -480 3850 -410
rect 1900 -490 3850 -480
rect 1790 -500 1900 -490
rect 3960 -490 3970 -410
rect 3850 -510 3960 -500
rect 770 -700 880 -690
rect 2830 -700 2940 -690
rect 760 -790 770 -710
rect 1280 -710 1392 -700
rect 2940 -710 2942 -700
rect 880 -790 1280 -710
rect 760 -800 1280 -790
rect 1392 -800 2830 -710
rect 2942 -720 3460 -710
rect 2942 -800 3340 -720
rect 760 -810 3340 -800
rect 3450 -810 3460 -720
rect 3340 -820 3450 -810
<< via2 >>
rect 758 370 760 460
rect 760 370 870 460
rect 3340 380 3450 460
rect 3450 380 3452 460
rect 3340 370 3452 380
rect 1280 60 1392 150
rect 2830 60 2942 150
rect 760 -480 872 -390
rect 3340 -480 3452 -390
rect 1280 -800 1390 -710
rect 1390 -800 1392 -710
rect 2830 -790 2940 -710
rect 2940 -790 2942 -710
rect 2830 -800 2942 -790
<< metal3 >>
rect 750 465 880 470
rect 748 460 880 465
rect 748 370 758 460
rect 870 370 880 460
rect 748 365 880 370
rect 750 -385 880 365
rect 3330 465 3460 470
rect 3330 460 3462 465
rect 3330 370 3340 460
rect 3452 370 3462 460
rect 3330 365 3462 370
rect 1270 155 1400 160
rect 1270 150 1402 155
rect 1270 60 1280 150
rect 1392 60 1402 150
rect 1270 55 1402 60
rect 2820 150 2952 155
rect 2820 60 2830 150
rect 2942 60 2952 150
rect 2820 55 2952 60
rect 750 -390 882 -385
rect 750 -480 760 -390
rect 872 -480 882 -390
rect 750 -485 882 -480
rect 750 -490 880 -485
rect 1270 -705 1400 55
rect 2820 -705 2950 55
rect 3330 -385 3460 365
rect 3330 -390 3462 -385
rect 3330 -480 3340 -390
rect 3452 -480 3462 -390
rect 3330 -485 3462 -480
rect 3330 -490 3460 -485
rect 1270 -710 1402 -705
rect 1270 -800 1280 -710
rect 1392 -800 1402 -710
rect 1270 -805 1402 -800
rect 2820 -710 2952 -705
rect 2820 -800 2830 -710
rect 2942 -800 2952 -710
rect 2820 -805 2952 -800
rect 1270 -810 1400 -805
rect 2820 -810 2950 -805
use sky130_fd_pr__pfet_01v8_lvt_B64SAM *sky130_fd_pr__pfet_01v8_lvt_B64SAM_0
timestamp 1661909013
transform 1 0 2109 0 1 224
box -2129 -264 2129 298
use sky130_fd_pr__pfet_01v8_lvt_MBDTEX  sky130_fd_pr__pfet_01v8_lvt_MBDTEX_0
timestamp 1661909182
transform 1 0 2109 0 1 -562
box -2129 -298 2129 264
<< labels >>
flabel nwell 3820 648 3980 828 0 FreeSans 1600 0 0 0 A
flabel nwell 3320 648 3480 828 0 FreeSans 1600 0 0 0 B
flabel nwell 2800 648 2960 828 0 FreeSans 1600 0 0 0 B
flabel nwell 2280 648 2440 828 0 FreeSans 1600 0 0 0 A
flabel nwell 1760 648 1920 828 0 FreeSans 1600 0 0 0 A
flabel nwell 1260 648 1420 828 0 FreeSans 1600 0 0 0 B
flabel nwell 740 648 900 828 0 FreeSans 1600 0 0 0 B
flabel nwell 240 648 400 828 0 FreeSans 1600 0 0 0 A
flabel space 3820 -1160 3980 -980 0 FreeSans 1600 0 0 0 B
flabel space 3300 -1160 3460 -980 0 FreeSans 1600 0 0 0 A
flabel space 2780 -1160 2940 -980 0 FreeSans 1600 0 0 0 A
flabel space 2280 -1160 2440 -980 0 FreeSans 1600 0 0 0 B
flabel space 1760 -1160 1920 -980 0 FreeSans 1600 0 0 0 B
flabel space 1240 -1160 1400 -980 0 FreeSans 1600 0 0 0 A
flabel space 720 -1160 880 -980 0 FreeSans 1600 0 0 0 A
flabel space 220 -1160 380 -980 0 FreeSans 1600 0 0 0 B
<< end >>
