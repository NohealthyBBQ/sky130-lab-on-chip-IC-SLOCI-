magic
tech sky130A
timestamp 1662865246
<< locali >>
rect -8750 6930 -8740 6960
rect -8750 6020 -8740 6050
rect -8750 5180 -8740 5210
rect -8750 4270 -8740 4300
rect -8750 3230 -8740 3260
rect -8750 2320 -8740 2350
rect -8750 1480 -8740 1510
rect -8750 570 -8740 600
rect -8750 -470 -8740 -440
rect -8750 -1380 -8740 -1350
rect -8750 -2220 -8740 -2190
rect -8750 -3130 -8740 -3100
rect -8710 6930 17660 6960
rect -8710 6020 17660 6050
rect -8710 5180 17660 5210
rect -8710 4270 17660 4300
rect -8710 3230 100 3260
rect 8850 3230 17660 3260
rect -8710 2320 100 2350
rect 8850 2320 17660 2350
rect -8710 1480 100 1510
rect 8850 1480 17660 1510
rect -8710 570 100 600
rect 8850 570 17660 600
rect -8710 -470 17660 -440
rect -8710 -1380 17660 -1350
rect -8710 -2220 17660 -2190
rect -8710 -3130 17660 -3100
rect 17690 6020 17700 6050
rect 17690 5180 17700 5210
rect 17690 4270 17700 4300
rect 17690 3230 17700 3260
rect 17690 2320 17700 2350
rect 17690 1480 17700 1510
rect 17690 570 17700 600
rect 17690 -470 17700 -440
rect 17690 -1380 17700 -1350
rect 17690 -2220 17700 -2190
rect 17690 -3130 17700 -3100
<< viali >>
rect -8660 7410 17620 7440
rect -8740 -3600 -8710 7400
rect 17660 -3600 17690 7400
rect -8670 -3640 17610 -3610
<< metal1 >>
rect -8750 7440 17700 7450
rect -8750 7410 -8660 7440
rect 17620 7410 17700 7440
rect -8750 7400 17700 7410
rect -8750 -3600 -8740 7400
rect -8710 6510 -8700 7400
rect 17650 6510 17660 7400
rect -8710 6470 17660 6510
rect -8710 4750 -8700 6470
rect 17650 4750 17660 6470
rect -8710 4710 17660 4750
rect -8710 -890 -8700 4710
rect 150 2710 210 2870
rect 1030 2820 1090 2870
rect 1030 2760 1300 2820
rect 2140 2760 2400 2820
rect 3240 2760 3500 2820
rect 4340 2760 4600 2820
rect 5440 2760 5700 2820
rect 6540 2760 6800 2820
rect 7640 2760 7900 2820
rect 1030 2710 1090 2760
rect 370 960 420 1100
rect 830 970 880 1110
rect 1040 1010 1310 1060
rect 2130 1010 2400 1060
rect 3230 1010 3500 1060
rect 4340 1010 4610 1060
rect 5440 1010 5710 1060
rect 6530 1010 6800 1060
rect 7640 1010 7910 1060
rect 17650 -890 17660 4710
rect -8710 -930 17660 -890
rect -8710 -2650 -8700 -930
rect 17650 -2650 17660 -930
rect -8710 -2690 17660 -2650
rect -8710 -3600 -8700 -2690
rect 17650 -3600 17660 -2690
rect 17690 -3600 17700 7400
rect -8750 -3610 17700 -3600
rect -8750 -3640 -8670 -3610
rect 17610 -3640 17700 -3610
rect -8750 -3650 17700 -3640
use XM_output_mirr_combined  XM_output_mirr_combined_0
timestamp 1662815693
transform 1 0 0 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_1
timestamp 1662815693
transform 1 0 0 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_2
timestamp 1662815693
transform 1 0 0 0 1 -3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_3
timestamp 1662815693
transform 1 0 -8800 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_4
timestamp 1662815693
transform 1 0 -8800 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_5
timestamp 1662815693
transform 1 0 -8800 0 1 -3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_6
timestamp 1662815693
transform 1 0 8800 0 1 3700
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_7
timestamp 1662815693
transform 1 0 8800 0 1 0
box 0 0 8950 3800
use XM_output_mirr_combined  XM_output_mirr_combined_8
timestamp 1662815693
transform 1 0 8800 0 1 -3700
box 0 0 8950 3800
<< labels >>
flabel space 40 44 8913 3752 0 FreeSans 6400 0 0 0 inner_core
<< end >>
