magic
tech sky130A
magscale 1 2
timestamp 1662671450
<< error_s >>
rect 67417 20989 67452 21023
rect 67418 20970 67452 20989
rect 822 15750 1566 15752
rect 822 14954 1566 14956
rect 7798 14799 7833 14833
rect 7799 14780 7833 14799
rect 822 14158 1566 14160
rect 822 13362 1566 13364
rect 3738 12781 3773 12815
rect 3739 12762 3773 12781
rect 822 12566 1566 12568
rect 822 11770 1566 11772
rect 822 10974 1566 10976
rect 822 10178 1566 10180
rect 822 9382 1566 9384
rect 822 8586 1566 8588
rect 822 7790 1566 7792
rect 822 6994 1566 6996
rect 822 6198 1566 6200
rect 822 5402 1566 5404
rect 822 4606 1566 4608
rect 822 3810 1566 3812
rect 822 3014 1566 3016
rect 822 2218 1566 2220
rect 1521 1931 1566 1985
rect 2714 1967 2748 1985
rect 1541 1424 1566 1931
rect 822 1422 1566 1424
rect 1575 1897 1620 1931
rect 822 626 824 1370
rect 1541 626 1566 1370
rect 1575 626 1609 1897
rect 1575 592 1600 626
rect 2678 583 2748 1967
rect 2678 547 2731 583
rect 3219 530 3234 5020
rect 3253 530 3287 5074
rect 3253 496 3268 530
rect 3758 477 3773 12762
rect 3792 12728 3827 12762
rect 4277 12728 4312 12762
rect 3792 477 3826 12728
rect 4278 12709 4312 12728
rect 3792 443 3807 477
rect 4297 424 4312 12709
rect 4331 12675 4366 12709
rect 4331 424 4365 12675
rect 6520 2541 6555 2575
rect 7113 2558 7147 2576
rect 6521 2522 6555 2541
rect 4786 978 4887 1232
rect 5040 488 5141 978
rect 5623 901 5657 920
rect 6035 902 6069 920
rect 5612 866 5657 901
rect 4331 390 4346 424
rect 5632 361 5657 866
rect 5666 832 5711 866
rect 5666 361 5700 832
rect 5812 764 5870 770
rect 5812 730 5824 764
rect 5812 724 5870 730
rect 5812 454 5870 460
rect 5812 420 5824 454
rect 5812 414 5870 420
rect 5666 327 5691 361
rect 5999 318 6069 902
rect 5999 282 6052 318
rect 6540 265 6555 2522
rect 6574 2488 6609 2522
rect 6574 265 6608 2488
rect 6574 231 6589 265
rect 7077 212 7147 2558
rect 7077 176 7130 212
rect 7818 159 7833 14780
rect 7852 14746 7887 14780
rect 7852 159 7886 14746
rect 10752 14481 10787 14515
rect 10753 14462 10787 14481
rect 10067 696 10101 714
rect 9106 664 9164 670
rect 8538 601 8572 655
rect 8960 637 8994 655
rect 7852 125 7867 159
rect 8557 106 8572 601
rect 8591 567 8626 601
rect 8591 106 8625 567
rect 8737 499 8795 505
rect 8737 465 8749 499
rect 8737 459 8795 465
rect 8737 189 8795 195
rect 8737 155 8749 189
rect 8737 149 8795 155
rect 8591 72 8606 106
rect 8924 53 8994 637
rect 9106 630 9118 664
rect 9106 624 9164 630
rect 9844 558 9902 564
rect 9276 531 9310 549
rect 9698 531 9732 549
rect 9276 495 9346 531
rect 9293 461 9364 495
rect 9106 136 9164 142
rect 9106 102 9118 136
rect 9106 96 9164 102
rect 8924 17 8977 53
rect 9293 0 9363 461
rect 9475 393 9533 399
rect 9475 359 9487 393
rect 9475 353 9533 359
rect 9475 83 9533 89
rect 9475 49 9487 83
rect 9475 43 9533 49
rect 9293 -36 9346 0
rect 9662 -53 9732 531
rect 9844 524 9856 558
rect 9844 518 9902 524
rect 9844 30 9902 36
rect 9844 -4 9856 30
rect 9844 -10 9902 -4
rect 9662 -89 9715 -53
rect 10031 -106 10101 696
rect 10031 -142 10084 -106
rect 10772 -159 10787 14462
rect 10806 14428 10841 14462
rect 11491 14428 11526 14462
rect 10806 -159 10840 14428
rect 11492 14409 11526 14428
rect 10806 -193 10821 -159
rect 11511 -212 11526 14409
rect 11545 14375 11580 14409
rect 12230 14375 12265 14409
rect 11545 -212 11579 14375
rect 12231 14356 12265 14375
rect 11545 -246 11560 -212
rect 12250 -265 12265 14356
rect 12284 14322 12319 14356
rect 12284 -265 12318 14322
rect 17207 14269 17242 14303
rect 17208 14250 17242 14269
rect 12284 -299 12299 -265
rect 17227 -371 17242 14250
rect 17261 14216 17296 14250
rect 17261 -371 17295 14216
rect 60819 14163 60854 14197
rect 60820 14144 60854 14163
rect 17261 -405 17276 -371
rect 60839 -477 60854 14144
rect 60873 14110 60908 14144
rect 61558 14110 61593 14144
rect 60873 -477 60907 14110
rect 61559 14091 61593 14110
rect 60873 -511 60888 -477
rect 61578 -530 61593 14091
rect 61612 14057 61647 14091
rect 62297 14057 62332 14091
rect 61612 -530 61646 14057
rect 62298 14038 62332 14057
rect 61612 -564 61627 -530
rect 62317 -583 62332 14038
rect 62351 14004 62386 14038
rect 63036 14004 63071 14038
rect 62351 -583 62385 14004
rect 63037 13985 63071 14004
rect 62351 -617 62366 -583
rect 63056 -636 63071 13985
rect 63090 13951 63125 13985
rect 63775 13951 63810 13985
rect 63090 -636 63124 13951
rect 63776 13932 63810 13951
rect 63090 -670 63105 -636
rect 63795 -689 63810 13932
rect 63829 13898 63864 13932
rect 64514 13898 64549 13932
rect 63829 -689 63863 13898
rect 64515 13879 64549 13898
rect 63829 -723 63844 -689
rect 64534 -742 64549 13879
rect 64568 13845 64603 13879
rect 65253 13845 65288 13879
rect 64568 -742 64602 13845
rect 65254 13826 65288 13845
rect 64568 -776 64583 -742
rect 65273 -795 65288 13826
rect 65307 13792 65342 13826
rect 65307 -795 65341 13792
rect 65307 -829 65322 -795
rect 66012 -848 66027 13826
rect 66046 -848 66080 13880
rect 66046 -882 66061 -848
rect 67437 -901 67452 20970
rect 67471 20936 67506 20970
rect 68842 20936 68877 20970
rect 67471 -901 67505 20936
rect 68843 20917 68877 20936
rect 67471 -935 67486 -901
rect 68862 -954 68877 20917
rect 68896 20883 68931 20917
rect 70267 20883 70302 20917
rect 68896 -954 68930 20883
rect 70268 20864 70302 20883
rect 68896 -988 68911 -954
rect 70287 -1007 70302 20864
rect 70321 20830 70356 20864
rect 71692 20830 71727 20864
rect 70321 -1007 70355 20830
rect 71693 20811 71727 20830
rect 70321 -1041 70336 -1007
rect 71712 -1060 71727 20811
rect 71746 20777 71781 20811
rect 71746 -1060 71780 20777
rect 71746 -1094 71761 -1060
rect 73137 -1113 73152 20811
rect 73171 -1113 73205 20865
rect 73679 8383 73713 8437
rect 73171 -1147 73186 -1113
rect 73698 -1166 73713 8383
rect 73732 8349 73767 8383
rect 73732 -1166 73766 8349
rect 74240 1472 74274 1526
rect 73732 -1200 73747 -1166
rect 74259 -1219 74274 1472
rect 74293 1438 74328 1472
rect 74293 -1219 74327 1438
rect 74293 -1253 74308 -1219
rect 74820 -1272 74835 1472
rect 74854 -1272 74888 1526
rect 74854 -1306 74869 -1272
use sky130_fd_pr__cap_mim_m3_1_ZQCY8R  XC_porst
timestamp 1662671450
transform 1 0 14790 0 1 1746
box -1750 -2100 1749 2100
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM4
timestamp 1662671450
transform 1 0 7473 0 1 7496
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM5
timestamp 1662671450
transform 1 0 8212 0 1 7443
box -396 -7373 396 7373
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM8
timestamp 1662671450
transform 1 0 6834 0 1 1367
box -296 -1191 296 1191
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM11
timestamp 1662671450
transform 1 0 6295 0 1 1420
box -296 -1191 296 1191
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM15
timestamp 1662671450
transform 1 0 10427 0 1 7178
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM16
timestamp 1662671450
transform 1 0 11166 0 1 7125
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM17
timestamp 1662671450
transform 1 0 11905 0 1 7072
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM18
timestamp 1662671450
transform 1 0 12644 0 1 7019
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM19
timestamp 1662671450
transform 1 0 16882 0 1 6966
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM20
timestamp 1662671450
transform 1 0 17621 0 1 6913
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM21
timestamp 1662671450
transform 1 0 60494 0 1 6860
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM22
timestamp 1662671450
transform 1 0 61233 0 1 6807
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM23
timestamp 1662671450
transform 1 0 61972 0 1 6754
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM24
timestamp 1662671450
transform 1 0 62711 0 1 6701
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM25
timestamp 1662671450
transform 1 0 63450 0 1 6648
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM26
timestamp 1662671450
transform 1 0 64189 0 1 6595
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM27
timestamp 1662671450
transform 1 0 64928 0 1 6542
box -396 -7373 396 7373
use sky130_fd_pr__nfet_01v8_lvt_WTP99N  XM28
timestamp 1662671450
transform 1 0 65667 0 1 6489
box -396 -7373 396 7373
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir1
timestamp 1662671450
transform 1 0 4052 0 1 6593
box -296 -6205 296 6205
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir2
timestamp 1662671450
transform 1 0 4591 0 1 6540
box -296 -6205 296 6205
use sky130_fd_pr__pfet_01v8_lvt_PH459S  XMfeedback_mir
timestamp 1662671450
transform 1 0 3513 0 1 6646
box -296 -6205 296 6205
use sky130_fd_pr__nfet_01v8_648S5X  XMinv_n1
timestamp 1662671450
transform 1 0 9504 0 1 221
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XMinv_n
timestamp 1662671450
transform 1 0 8766 0 1 327
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XMinv_p1
timestamp 1662671450
transform 1 0 9873 0 1 277
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XMinv_p
timestamp 1662671450
transform 1 0 9135 0 1 383
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_lvt_AHZKRZ  XMota_bias_n
timestamp 1662671450
transform 1 0 2135 0 1 1257
box -596 -710 596 710
use sky130_fd_pr__pfet_01v8_lvt_AH4MH9  XMota_bias_p
timestamp 1662671450
transform 1 0 2974 0 1 2775
box -296 -2281 296 2281
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XMpdn
timestamp 1662671450
transform 1 0 5841 0 1 592
box -211 -310 211 310
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 0 796 0 33 796
timestamp 1657128861
transform 1 0 796 0 1 600
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
timestamp 1657128861
transform 1 0 0 0 1 600
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1657128861
transform 1 0 4887 0 1 335
box 0 0 796 796
use sky130_fd_pr__res_high_po_1p41_LKUZST  XR3
timestamp 1662671450
transform 1 0 74564 0 1 100
box -307 -1408 307 1408
use sky130_fd_pr__res_high_po_1p41_S8KB58  XR4
timestamp 1662671450
transform 1 0 74003 0 1 3582
box -307 -4837 307 4837
use sky130_fd_pr__res_high_po_1p41_6AVB5Q  XR_porst
timestamp 1662671450
transform 1 0 75125 0 1 837
box -307 -2198 307 2198
use sky130_fd_pr__res_high_po_1p41_7S2UWS  XRref_high
timestamp 1662671450
transform 1 0 73442 0 1 14746
box -307 -15948 307 15948
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh1
timestamp 1662671450
transform 1 0 68174 0 1 10008
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh2
timestamp 1662671450
transform 1 0 69599 0 1 9955
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh3
timestamp 1662671450
transform 1 0 71024 0 1 9902
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh4
timestamp 1662671450
transform 1 0 72449 0 1 9849
box -739 -10998 739 10998
use sky130_fd_pr__res_xhigh_po_5p73_AUAUMD  XRref_xhigh
timestamp 1662671450
transform 1 0 66749 0 1 10061
box -739 -10998 739 10998
<< end >>
