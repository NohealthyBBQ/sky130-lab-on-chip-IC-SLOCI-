magic
tech sky130A
magscale 1 2
timestamp 1662674005
<< nwell >>
rect -162 -100 2374 2674
<< metal1 >>
rect 790 2440 800 2500
rect 860 2440 870 2500
rect 1830 2440 1840 2500
rect 1900 2440 1910 2500
rect 290 2300 300 2360
rect 360 2300 370 2360
rect 1310 2300 1320 2360
rect 1380 2300 1390 2360
rect 98 2202 2096 2250
rect 790 2060 800 2120
rect 860 2060 870 2120
rect 1830 2060 1840 2120
rect 1900 2060 1910 2120
rect 290 1920 300 1980
rect 360 1920 370 1980
rect 1310 1920 1320 1980
rect 1380 1920 1390 1980
rect 98 1838 2096 1884
rect 790 1700 800 1760
rect 860 1700 870 1760
rect 1830 1700 1840 1760
rect 1900 1700 1910 1760
rect 290 1560 300 1620
rect 360 1560 370 1620
rect 1310 1560 1320 1620
rect 1380 1560 1390 1620
rect 98 1472 2096 1520
rect 810 1340 820 1400
rect 880 1340 890 1400
rect 1830 1340 1840 1400
rect 1900 1340 1910 1400
rect 290 1200 300 1260
rect 360 1200 370 1260
rect 1330 1200 1340 1260
rect 1400 1200 1410 1260
rect 98 1108 2096 1154
rect 790 980 800 1040
rect 860 980 870 1040
rect 1830 980 1840 1040
rect 1900 980 1910 1040
rect 290 840 300 900
rect 360 840 370 900
rect 1310 840 1320 900
rect 1380 840 1390 900
rect 98 742 2096 790
rect 790 600 800 660
rect 860 600 870 660
rect 1830 600 1840 660
rect 1900 600 1910 660
rect 290 460 300 520
rect 360 460 370 520
rect 1310 460 1320 520
rect 1380 460 1390 520
rect 98 378 2096 424
rect 790 240 800 300
rect 860 240 870 300
rect 1830 240 1840 300
rect 1900 240 1910 300
rect 290 100 300 160
rect 360 100 370 160
rect 1310 100 1320 160
rect 1380 100 1390 160
rect 98 12 2096 60
<< via1 >>
rect 800 2440 860 2500
rect 1840 2440 1900 2500
rect 300 2300 360 2360
rect 1320 2300 1380 2360
rect 800 2060 860 2120
rect 1840 2060 1900 2120
rect 300 1920 360 1980
rect 1320 1920 1380 1980
rect 800 1700 860 1760
rect 1840 1700 1900 1760
rect 300 1560 360 1620
rect 1320 1560 1380 1620
rect 820 1340 880 1400
rect 1840 1340 1900 1400
rect 300 1200 360 1260
rect 1340 1200 1400 1260
rect 800 980 860 1040
rect 1840 980 1900 1040
rect 300 840 360 900
rect 1320 840 1380 900
rect 800 600 860 660
rect 1840 600 1900 660
rect 300 460 360 520
rect 1320 460 1380 520
rect 800 240 860 300
rect 1840 240 1900 300
rect 300 100 360 160
rect 1320 100 1380 160
<< metal2 >>
rect 800 2510 1880 2520
rect 800 2500 1900 2510
rect 860 2480 1840 2500
rect 800 2430 860 2440
rect 1840 2430 1900 2440
rect 300 2360 360 2370
rect 1320 2360 1380 2370
rect 360 2300 1320 2320
rect 300 2280 1380 2300
rect 800 2120 1900 2140
rect 860 2100 1840 2120
rect 800 2050 860 2060
rect 1840 2050 1900 2060
rect 300 1980 360 1990
rect 1320 1980 1380 1990
rect 360 1920 1320 1940
rect 300 1900 1380 1920
rect 800 1760 1900 1780
rect 860 1740 1840 1760
rect 800 1690 860 1700
rect 1840 1690 1900 1700
rect 300 1620 360 1630
rect 1320 1620 1380 1630
rect 360 1560 1320 1580
rect 300 1540 1380 1560
rect 820 1400 1900 1420
rect 880 1380 1840 1400
rect 820 1330 880 1340
rect 1840 1330 1900 1340
rect 300 1260 360 1270
rect 1340 1260 1400 1270
rect 360 1200 1340 1220
rect 300 1180 1400 1200
rect 800 1040 1900 1060
rect 860 1020 1840 1040
rect 800 970 860 980
rect 1840 970 1900 980
rect 300 900 360 910
rect 1320 900 1380 910
rect 360 840 1320 860
rect 300 820 1380 840
rect 800 660 1900 680
rect 860 640 1840 660
rect 800 590 860 600
rect 1840 590 1900 600
rect 300 520 360 530
rect 1320 520 1380 530
rect 360 460 1320 480
rect 300 440 1380 460
rect 800 300 1900 320
rect 860 280 1840 300
rect 800 230 860 240
rect 1840 230 1900 240
rect 300 160 360 170
rect 1320 160 1380 170
rect 360 100 1320 120
rect 300 80 1380 100
<< metal3 >>
rect 40 100 100 2500
rect 560 100 620 2500
rect 1060 100 1120 2500
rect 1580 100 1640 2500
rect 2100 100 2160 2500
use sky130_fd_pr__pfet_01v8_lvt_8URDWJ  sky130_fd_pr__pfet_01v8_lvt_8URDWJ_0
timestamp 1662671833
transform 1 0 1097 0 1 1260
box -1097 -1260 1097 1292
<< labels >>
flabel nwell 300 2540 360 2620 0 FreeSans 800 0 0 0 A
flabel nwell 1340 2540 1400 2620 0 FreeSans 800 0 0 0 A
flabel nwell 820 2160 880 2240 0 FreeSans 800 0 0 0 A
flabel nwell 1840 2140 1900 2220 0 FreeSans 800 0 0 0 A
flabel nwell 280 1780 340 1860 0 FreeSans 800 0 0 0 A
flabel nwell 1340 1800 1400 1880 0 FreeSans 800 0 0 0 A
flabel nwell 820 1400 880 1480 0 FreeSans 800 0 0 0 A
flabel nwell 1840 1400 1900 1480 0 FreeSans 800 0 0 0 A
flabel nwell 300 1040 360 1120 0 FreeSans 800 0 0 0 A
flabel nwell 1340 1060 1400 1140 0 FreeSans 800 0 0 0 A
flabel nwell 780 680 840 760 0 FreeSans 800 0 0 0 A
flabel nwell 1860 680 1920 760 0 FreeSans 800 0 0 0 A
flabel nwell 280 300 340 380 0 FreeSans 800 0 0 0 A
flabel nwell 1320 300 1380 380 0 FreeSans 800 0 0 0 A
flabel nwell 820 2520 880 2600 0 FreeSans 800 0 0 0 B
flabel nwell 1840 2520 1900 2600 0 FreeSans 800 0 0 0 B
flabel nwell 300 2140 360 2220 0 FreeSans 800 0 0 0 B
flabel nwell 1340 2140 1400 2220 0 FreeSans 800 0 0 0 B
flabel nwell 820 1780 880 1860 0 FreeSans 800 0 0 0 B
flabel nwell 1860 1780 1920 1860 0 FreeSans 800 0 0 0 B
flabel nwell 280 1400 340 1480 0 FreeSans 800 0 0 0 B
flabel nwell 1340 1420 1400 1500 0 FreeSans 800 0 0 0 B
flabel nwell 820 1060 880 1140 0 FreeSans 800 0 0 0 B
flabel nwell 1840 1060 1900 1140 0 FreeSans 800 0 0 0 B
flabel nwell 300 700 360 780 0 FreeSans 800 0 0 0 B
flabel nwell 1340 680 1400 760 0 FreeSans 800 0 0 0 B
flabel nwell 820 320 880 400 0 FreeSans 800 0 0 0 B
flabel nwell 1840 320 1900 400 0 FreeSans 800 0 0 0 B
<< end >>
