magic
tech sky130A
magscale 1 2
timestamp 1662136735
<< pwell >>
rect -400 -1400 1600 1700
<< psubdiff >>
rect -320 1540 1480 1560
rect -320 1500 -220 1540
rect 0 1500 240 1540
rect 460 1500 700 1540
rect 920 1500 1160 1540
rect 1380 1500 1480 1540
rect -320 1480 1480 1500
rect -320 1200 -240 1480
rect -320 980 -300 1200
rect -260 980 -240 1200
rect -320 720 -240 980
rect -320 500 -300 720
rect -260 500 -240 720
rect -320 180 -240 500
rect 1400 1200 1480 1480
rect 1400 980 1420 1200
rect 1460 980 1480 1200
rect 1400 720 1480 980
rect 1400 500 1420 720
rect 1460 500 1480 720
rect 1400 180 1480 500
rect -320 160 1480 180
rect -320 120 -220 160
rect 0 120 240 160
rect 460 120 700 160
rect 920 120 1160 160
rect 1380 120 1480 160
rect -320 100 1480 120
rect -320 -140 -240 100
rect -320 -360 -300 -140
rect -260 -360 -240 -140
rect -320 -700 -240 -360
rect -320 -920 -300 -700
rect -260 -920 -240 -700
rect -320 -1200 -240 -920
rect 1400 -140 1480 100
rect 1400 -360 1420 -140
rect 1460 -360 1480 -140
rect 1400 -700 1480 -360
rect 1400 -920 1420 -700
rect 1460 -920 1480 -700
rect 1400 -1200 1480 -920
rect -320 -1220 1480 -1200
rect -320 -1260 -220 -1220
rect 0 -1260 240 -1220
rect 460 -1260 700 -1220
rect 920 -1260 1160 -1220
rect 1380 -1260 1480 -1220
rect -320 -1280 1480 -1260
<< psubdiffcont >>
rect -220 1500 0 1540
rect 240 1500 460 1540
rect 700 1500 920 1540
rect 1160 1500 1380 1540
rect -300 980 -260 1200
rect -300 500 -260 720
rect 1420 980 1460 1200
rect 1420 500 1460 720
rect -220 120 0 160
rect 240 120 460 160
rect 700 120 920 160
rect 1160 120 1380 160
rect -300 -360 -260 -140
rect -300 -920 -260 -700
rect 1420 -360 1460 -140
rect 1420 -920 1460 -700
rect -220 -1260 0 -1220
rect 240 -1260 460 -1220
rect 700 -1260 920 -1220
rect 1160 -1260 1380 -1220
<< locali >>
rect -320 1540 1480 1560
rect -320 1500 -220 1540
rect 0 1500 240 1540
rect 460 1500 700 1540
rect 920 1500 1160 1540
rect 1380 1500 1480 1540
rect -320 1480 1480 1500
rect -320 1200 -240 1480
rect -320 980 -300 1200
rect -260 980 -240 1200
rect -320 720 -240 980
rect -320 500 -300 720
rect -260 500 -240 720
rect -320 180 -240 500
rect 1400 1200 1480 1480
rect 1400 980 1420 1200
rect 1460 980 1480 1200
rect 1400 720 1480 980
rect 1400 500 1420 720
rect 1460 500 1480 720
rect 1400 180 1480 500
rect -320 160 1480 180
rect -320 120 -220 160
rect 0 120 240 160
rect 460 120 700 160
rect 920 120 1160 160
rect 1380 120 1480 160
rect -320 100 1480 120
rect -320 -140 -240 100
rect -320 -360 -300 -140
rect -260 -360 -240 -140
rect -320 -700 -240 -360
rect -320 -920 -300 -700
rect -260 -920 -240 -700
rect -320 -1200 -240 -920
rect 1400 -140 1480 100
rect 1400 -360 1420 -140
rect 1460 -360 1480 -140
rect 1400 -700 1480 -360
rect 1400 -920 1420 -700
rect 1460 -920 1480 -700
rect 1400 -1200 1480 -920
rect -320 -1220 1480 -1200
rect -320 -1260 -220 -1220
rect 0 -1260 240 -1220
rect 460 -1260 700 -1220
rect 920 -1260 1160 -1220
rect 1380 -1260 1480 -1220
rect -320 -1280 1480 -1260
<< viali >>
rect -220 1500 0 1540
rect 240 1500 460 1540
rect 700 1500 920 1540
rect 1160 1500 1380 1540
rect -300 980 -260 1200
rect -300 500 -260 720
rect 1420 980 1460 1200
rect 1420 500 1460 720
rect -300 -360 -260 -140
rect -300 -920 -260 -700
rect 1420 -360 1460 -140
rect 1420 -920 1460 -700
rect -220 -1260 0 -1220
rect 240 -1260 460 -1220
rect 700 -1260 920 -1220
rect 1160 -1260 1380 -1220
<< metal1 >>
rect -320 1540 1480 1560
rect -320 1500 -220 1540
rect 0 1500 240 1540
rect 460 1500 700 1540
rect 920 1500 1160 1540
rect 1380 1500 1480 1540
rect -320 1480 1480 1500
rect -320 1200 -240 1480
rect 30 1280 40 1340
rect 100 1280 110 1340
rect 304 1326 350 1480
rect 820 1326 866 1480
rect 1060 1280 1070 1340
rect 1130 1280 1140 1340
rect -320 980 -300 1200
rect -260 980 -240 1200
rect -320 720 -240 980
rect -320 500 -300 720
rect -260 500 -240 720
rect -320 -140 -240 500
rect 1400 1200 1480 1480
rect 1400 980 1420 1200
rect 1460 980 1480 1200
rect 1400 720 1480 980
rect 1400 500 1420 720
rect 1460 500 1480 720
rect 544 438 554 498
rect 614 438 624 498
rect 160 260 240 400
rect 160 200 170 260
rect 230 200 240 260
rect 430 80 510 400
rect 551 360 619 406
rect 930 260 1010 400
rect 160 20 170 80
rect 230 20 240 80
rect 430 20 440 80
rect 500 20 510 80
rect 660 200 670 260
rect 730 200 740 260
rect 930 200 940 260
rect 1000 200 1010 260
rect 160 -120 240 20
rect 551 -122 619 -76
rect 660 -120 740 200
rect 930 20 940 80
rect 1000 20 1010 80
rect 930 -120 1010 20
rect -320 -360 -300 -140
rect -260 -360 -240 -140
rect 1400 -140 1480 500
rect 545 -214 555 -154
rect 615 -214 625 -154
rect -320 -700 -240 -360
rect -320 -920 -300 -700
rect -260 -920 -240 -700
rect -320 -1200 -240 -920
rect 1400 -360 1420 -140
rect 1460 -360 1480 -140
rect 1400 -700 1480 -360
rect 1400 -920 1420 -700
rect 1460 -920 1480 -700
rect 30 -1060 40 -1000
rect 100 -1060 110 -1000
rect 304 -1200 350 -1042
rect 820 -1200 866 -1042
rect 1060 -1060 1070 -1000
rect 1130 -1060 1140 -1000
rect 1400 -1200 1480 -920
rect -320 -1220 1480 -1200
rect -320 -1260 -220 -1220
rect 0 -1260 240 -1220
rect 460 -1260 700 -1220
rect 920 -1260 1160 -1220
rect 1380 -1260 1480 -1220
rect -320 -1280 1480 -1260
<< via1 >>
rect 40 1280 100 1340
rect 1070 1280 1130 1340
rect 554 438 614 498
rect 170 200 230 260
rect 170 20 230 80
rect 440 20 500 80
rect 670 200 730 260
rect 940 200 1000 260
rect 940 20 1000 80
rect 555 -214 615 -154
rect 40 -1060 100 -1000
rect 1070 -1060 1130 -1000
<< metal2 >>
rect 40 1340 1266 1350
rect 100 1280 1070 1340
rect 1130 1280 1266 1340
rect 40 1270 1266 1280
rect -98 498 614 508
rect -98 438 554 498
rect -98 428 614 438
rect -98 -990 -30 428
rect 170 260 1000 270
rect 230 200 670 260
rect 730 200 940 260
rect 170 190 1000 200
rect 170 80 1000 90
rect 230 20 440 80
rect 500 20 940 80
rect 170 10 1000 20
rect 1198 -144 1266 1270
rect 554 -154 1266 -144
rect 554 -214 555 -154
rect 615 -214 1266 -154
rect 554 -224 1266 -214
rect -98 -1000 1130 -990
rect -98 -1060 40 -1000
rect 100 -1060 1070 -1000
rect -98 -1070 1130 -1060
use sky130_fd_pr__nfet_01v8_lvt_A5VCMN  sky130_fd_pr__nfet_01v8_lvt_A5VCMN_0
timestamp 1662090071
transform 1 0 585 0 1 -573
box -545 -507 545 507
use sky130_fd_pr__nfet_01v8_lvt_E96B6C  sky130_fd_pr__nfet_01v8_lvt_E96B6C_0
timestamp 1662090071
transform 1 0 585 0 1 857
box -545 -507 545 507
<< labels >>
flabel space 116 1692 300 1816 0 FreeSans 1280 0 0 0 A
flabel space 360 1688 544 1812 0 FreeSans 1280 0 0 0 B
flabel space 624 1696 808 1820 0 FreeSans 1280 0 0 0 B
flabel space 886 1686 1070 1810 0 FreeSans 1280 0 0 0 A
flabel space 98 -1638 282 -1514 0 FreeSans 1280 0 0 0 B
flabel space 388 -1626 572 -1502 0 FreeSans 1280 0 0 0 A
flabel space 654 -1638 838 -1514 0 FreeSans 1280 0 0 0 A
flabel space 890 -1642 1074 -1518 0 FreeSans 1280 0 0 0 B
flabel pwell 1320 200 1400 260 0 FreeSans 480 0 0 0 A
flabel pwell 1320 20 1400 80 0 FreeSans 480 0 0 0 B
<< end >>
