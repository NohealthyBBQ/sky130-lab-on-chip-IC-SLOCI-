magic
tech sky130A
magscale 1 2
timestamp 1662767476
<< metal1 >>
rect 62 -98 1828 56
rect 62 -3610 1828 -3456
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_0
timestamp 1662766393
transform 1 0 945 0 1 -899
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_1
timestamp 1662766393
transform 1 0 945 0 1 -4411
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_0
timestamp 1662766393
transform 1 0 945 0 1 857
box -945 -857 945 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_1
timestamp 1662766393
transform 1 0 945 0 1 -2655
box -945 -857 945 857
<< end >>
