magic
tech sky130A
magscale 1 2
timestamp 1662665204
<< locali >>
rect 4525 -40 4560 105
rect 5040 -40 5075 105
rect 4525 -660 4560 -515
rect 5040 -655 5075 -510
rect 4525 -1155 4560 -1045
rect 4250 -1190 4560 -1155
rect 5040 -1185 5075 -1040
rect 4250 -1300 4560 -1285
rect 4250 -1340 4335 -1300
rect 4475 -1340 4560 -1300
rect 4250 -1355 4560 -1340
rect 4250 -1505 4560 -1470
<< viali >>
rect 4335 -1340 4475 -1300
<< metal1 >>
rect 3300 860 5110 920
rect 4610 300 4670 860
rect 4700 810 4780 820
rect 4700 750 4710 810
rect 4770 800 4780 810
rect 4770 750 4900 800
rect 4700 740 4780 750
rect 4820 710 4900 720
rect 4820 700 4830 710
rect 4700 650 4830 700
rect 4890 650 4900 710
rect 4820 640 4900 650
rect 4700 610 4780 620
rect 4700 550 4710 610
rect 4770 600 4780 610
rect 4770 560 4900 600
rect 4770 550 4780 560
rect 4700 540 4780 550
rect 4820 510 4900 520
rect 4700 460 4830 510
rect 4820 450 4830 460
rect 4890 450 4900 510
rect 4820 440 4900 450
rect 4700 420 4780 430
rect 4700 360 4710 420
rect 4770 410 4780 420
rect 4770 370 4900 410
rect 4770 360 4780 370
rect 4700 350 4780 360
rect 4820 320 4900 330
rect 4700 270 4830 320
rect 4820 260 4830 270
rect 4890 260 4900 320
rect 4820 250 4900 260
rect 4700 220 4780 230
rect 4700 160 4710 220
rect 4770 170 4900 220
rect 4930 210 4990 860
rect 4770 160 4780 170
rect 4700 150 4780 160
rect 3300 -50 5110 10
rect 4610 -410 4670 -50
rect 4700 -110 4780 -100
rect 4700 -170 4710 -110
rect 4770 -170 4780 -110
rect 4700 -180 4780 -170
rect 4820 -200 4900 -190
rect 4820 -260 4830 -200
rect 4890 -260 4900 -200
rect 4820 -270 4900 -260
rect 4700 -300 4780 -290
rect 4700 -360 4710 -300
rect 4770 -360 4780 -300
rect 4930 -310 4990 -50
rect 4700 -370 4780 -360
rect 4820 -390 4900 -380
rect 4820 -450 4830 -390
rect 4890 -450 4900 -390
rect 4820 -460 4900 -450
rect 3300 -640 5110 -580
rect 4610 -670 4990 -640
rect 4610 -830 4670 -670
rect 4700 -720 4780 -710
rect 4700 -780 4710 -720
rect 4770 -780 4780 -720
rect 4700 -790 4780 -780
rect 4820 -820 4900 -810
rect 4820 -880 4830 -820
rect 4890 -880 4900 -820
rect 4820 -890 4900 -880
rect 4700 -910 4780 -900
rect 4700 -970 4710 -910
rect 4770 -970 4780 -910
rect 4930 -930 4990 -670
rect 4700 -980 4780 -970
rect 3300 -1180 5110 -1120
rect 3910 -1250 3990 -1240
rect 3820 -1360 3880 -1290
rect 3910 -1310 3920 -1250
rect 3980 -1262 3990 -1250
rect 4700 -1250 4780 -1240
rect 3980 -1308 4110 -1262
rect 4320 -1290 4490 -1285
rect 3980 -1310 3990 -1308
rect 3910 -1320 3990 -1310
rect 4030 -1350 4110 -1340
rect 3910 -1396 4040 -1350
rect 4030 -1410 4040 -1396
rect 4100 -1410 4110 -1350
rect 4030 -1420 4110 -1410
rect 4140 -1480 4200 -1290
rect 4320 -1350 4335 -1290
rect 4475 -1350 4490 -1290
rect 4320 -1355 4490 -1350
rect 4610 -1360 4670 -1290
rect 4700 -1310 4710 -1250
rect 4770 -1310 4780 -1250
rect 4700 -1320 4780 -1310
rect 4820 -1350 4900 -1340
rect 4820 -1410 4830 -1350
rect 4890 -1410 4900 -1350
rect 4930 -1360 4990 -1180
rect 4820 -1420 4900 -1410
rect 3300 -1540 5110 -1480
<< via1 >>
rect 4710 750 4770 810
rect 4830 650 4890 710
rect 4710 550 4770 610
rect 4830 450 4890 510
rect 4710 360 4770 420
rect 4830 260 4890 320
rect 4710 160 4770 220
rect 4710 -170 4770 -110
rect 4830 -260 4890 -200
rect 4710 -360 4770 -300
rect 4830 -450 4890 -390
rect 4710 -780 4770 -720
rect 4830 -880 4890 -820
rect 4710 -970 4770 -910
rect 3920 -1310 3980 -1250
rect 4040 -1410 4100 -1350
rect 4335 -1300 4475 -1290
rect 4335 -1340 4475 -1300
rect 4335 -1350 4475 -1340
rect 4710 -1310 4770 -1250
rect 4830 -1410 4890 -1350
<< metal2 >>
rect 4520 810 4780 920
rect 4950 910 5110 920
rect 4520 750 4710 810
rect 4770 750 4780 810
rect 4520 610 4780 750
rect 4520 550 4710 610
rect 4770 550 4780 610
rect 4520 420 4780 550
rect 4520 360 4710 420
rect 4770 360 4780 420
rect 4520 220 4780 360
rect 4520 160 4710 220
rect 4770 160 4780 220
rect 4520 -110 4780 160
rect 4820 710 4980 910
rect 4820 650 4830 710
rect 4890 650 4980 710
rect 4820 510 4980 650
rect 4820 450 4830 510
rect 4890 450 4980 510
rect 4820 320 4980 450
rect 4820 260 4830 320
rect 4890 260 4980 320
rect 4820 90 4980 260
rect 5080 90 5110 910
rect 4820 60 5110 90
rect 4520 -170 4710 -110
rect 4770 -170 4780 -110
rect 4520 -300 4780 -170
rect 4520 -360 4710 -300
rect 4770 -360 4780 -300
rect 4520 -720 4780 -360
rect 4820 -30 5110 10
rect 4820 -200 4980 -30
rect 4820 -260 4830 -200
rect 4890 -260 4980 -200
rect 4820 -390 4980 -260
rect 4820 -450 4830 -390
rect 4890 -450 4980 -390
rect 4820 -530 4980 -450
rect 5080 -530 5110 -30
rect 4820 -550 5110 -530
rect 4820 -560 5080 -550
rect 4520 -780 4710 -720
rect 4770 -780 4780 -720
rect 4520 -910 4780 -780
rect 4520 -970 4710 -910
rect 4770 -970 4780 -910
rect 4520 -1150 4780 -970
rect 4820 -650 5110 -610
rect 4820 -820 4980 -650
rect 4820 -880 4830 -820
rect 4890 -880 4980 -820
rect 4820 -1030 4980 -880
rect 5080 -1030 5110 -650
rect 4820 -1060 5110 -1030
rect 4820 -1070 5080 -1060
rect 3730 -1180 3990 -1150
rect 3730 -1470 3760 -1180
rect 3880 -1250 3990 -1180
rect 3880 -1310 3920 -1250
rect 3980 -1310 3990 -1250
rect 3880 -1470 3990 -1310
rect 3730 -1510 3990 -1470
rect 4030 -1250 4780 -1150
rect 4030 -1290 4710 -1250
rect 4030 -1350 4335 -1290
rect 4475 -1310 4710 -1290
rect 4770 -1310 4780 -1250
rect 4475 -1350 4780 -1310
rect 4030 -1410 4040 -1350
rect 4100 -1410 4780 -1350
rect 4030 -1510 4780 -1410
rect 4820 -1180 5080 -1150
rect 4820 -1350 4950 -1180
rect 4820 -1410 4830 -1350
rect 4890 -1410 4950 -1350
rect 4820 -1480 4950 -1410
rect 5050 -1480 5080 -1180
rect 4820 -1510 5080 -1480
<< via2 >>
rect 4980 90 5080 910
rect 4980 -530 5080 -30
rect 4980 -1030 5080 -650
rect 3760 -1470 3880 -1180
rect 4950 -1480 5050 -1180
<< metal3 >>
rect 4950 910 5110 920
rect 4950 90 4980 910
rect 5080 90 5110 910
rect 4950 60 5110 90
rect 4950 -30 5110 0
rect 4950 -530 4980 -30
rect 5080 -530 5110 -30
rect 4950 -550 5110 -530
rect 4950 -650 5110 -630
rect 4950 -1030 4980 -650
rect 5080 -1030 5110 -650
rect 4950 -1060 5110 -1030
rect 3730 -1180 3900 -1150
rect 3730 -1470 3760 -1180
rect 3880 -1470 3900 -1180
rect 3730 -1510 3900 -1470
rect 4920 -1180 5080 -1150
rect 4920 -1480 4950 -1180
rect 5050 -1480 5080 -1180
rect 4920 -1510 5080 -1480
<< via3 >>
rect 4980 90 5080 910
rect 4980 -530 5080 -30
rect 4980 -1030 5080 -650
rect 3760 -1470 3880 -1180
rect 4950 -1480 5050 -1180
<< metal4 >>
rect 4370 2260 4890 2540
rect 3730 -1180 4090 -500
rect 4510 -630 4670 1930
rect 4730 0 4890 2260
rect 4950 910 5110 4368
rect 4950 90 4980 910
rect 5080 90 5110 910
rect 4950 60 5110 90
rect 4730 -30 5110 0
rect 4730 -530 4980 -30
rect 5080 -530 5110 -30
rect 4730 -560 5110 -530
rect 4510 -650 5110 -630
rect 4510 -1030 4980 -650
rect 5080 -1030 5110 -650
rect 4510 -1060 5110 -1030
rect 4510 -1070 5080 -1060
rect 3730 -1470 3760 -1180
rect 3880 -1470 4090 -1180
rect 3730 -1510 4090 -1470
rect 4760 -1180 5080 -1150
rect 4760 -1480 4810 -1180
rect 5050 -1480 5080 -1180
rect 4760 -1510 5080 -1480
<< via4 >>
rect 4810 -1480 4950 -1180
rect 4950 -1480 5050 -1180
<< metal5 >>
rect 3380 3710 4990 4830
rect 3380 3700 4930 3710
rect 3380 1430 3970 3700
rect 3380 -420 3780 1430
rect 4280 400 5080 1000
rect 4760 -1180 5080 400
rect 4760 -1480 4810 -1180
rect 5050 -1480 5080 -1180
rect 4760 -1510 5080 -1480
use sky130_fd_pr__cap_mim_m3_2_WCTBV5  XC1
timestamp 1660521579
transform 1 0 3851 0 1 701
box -551 -301 573 301
use sky130_fd_pr__cap_mim_m3_2_WCTZRP  XC2
timestamp 1660420676
transform 1 0 3951 0 1 1631
box -651 -301 673 301
use sky130_fd_pr__cap_mim_m3_2_3ZFDVT  XC3
timestamp 1660420676
transform 1 0 3951 0 1 2761
box -651 -501 673 501
use sky130_fd_pr__cap_mim_m3_2_VCH7EQ  XC4
timestamp 1660420676
transform 0 1 4611 1 0 4541
box -951 -501 973 501
use sky130_fd_pr__cap_mim_m3_2_FJFAMD  XC6
timestamp 1660420676
transform 1 0 3851 0 1 -229
box -551 -301 573 301
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1 backup/1.7_10G
timestamp 1662404926
transform 0 1 4010 -1 0 -1329
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM2
timestamp 1662404926
transform 0 1 4800 -1 0 -1329
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM3
timestamp 1660420676
transform 0 -1 4800 1 0 -847
box -263 -310 263 310
use sky130_fd_pr__nfet_01v8_lvt_BX7S53  XM4
timestamp 1660420676
transform 0 1 4800 -1 0 -279
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_lvt_B6HS5D  XM5
timestamp 1660420676
transform 0 1 4800 -1 0 485
box -455 -310 455 310
<< labels >>
rlabel metal2 4100 -1510 4710 -1150 1 GND
rlabel metal5 3380 3700 4930 4830 1 IN
rlabel metal1 3300 -1540 5110 -1480 1 ctrll1
rlabel metal1 3300 -1180 5110 -1120 1 ctrll2
rlabel metal1 3300 -640 5110 -580 1 ctrll3
rlabel metal1 3300 -50 5110 10 1 ctrll4
rlabel metal1 3300 860 5110 920 1 ctrll5
<< end >>
