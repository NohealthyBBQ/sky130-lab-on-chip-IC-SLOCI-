magic
tech sky130A
magscale 1 2
timestamp 1662990520
<< locali >>
rect 3988 -59524 4946 -59486
rect 5164 -59618 5202 -59504
rect 5578 -59612 5616 -59498
rect 6008 -59606 6046 -59492
rect 6428 -59608 6466 -59494
rect 6844 -59608 6882 -59494
rect 7262 -59608 7300 -59494
rect 7680 -59608 7718 -59494
rect 8096 -59608 8134 -59494
rect 8514 -59608 8552 -59494
rect 8932 -59608 8970 -59494
rect 9350 -59608 9388 -59494
rect 9766 -59608 9804 -59494
rect 10184 -59608 10222 -59494
rect 10602 -59608 10640 -59494
rect 11018 -59608 11056 -59494
rect 11436 -59608 11474 -59494
rect 11854 -59608 11892 -59494
rect 12270 -59608 12308 -59494
rect 12688 -59608 12726 -59494
rect 13106 -59608 13144 -59494
rect 13524 -59608 13562 -59494
rect 13940 -59608 13978 -59494
rect 14358 -59608 14396 -59494
rect 14776 -59608 14814 -59494
rect 15192 -59608 15230 -59494
rect 15610 -59608 15648 -59494
rect 16028 -59608 16066 -59494
rect 16444 -59608 16482 -59494
rect 9190 -59816 9424 -59814
rect 9190 -59936 9444 -59816
rect 9210 -59938 9444 -59936
<< viali >>
rect 3660 -59522 3724 -59456
<< metal1 >>
rect 20608 9410 23560 9440
rect 48 8820 288 8850
rect -268 -5380 -258 -5328
rect -206 -5380 -196 -5328
rect -686 -19582 -676 -19530
rect -624 -19582 -614 -19530
rect -1094 -33752 -1084 -33700
rect -1032 -33752 -1022 -33700
rect -1090 -49700 -1060 -33752
rect -678 -35496 -648 -19582
rect -258 -21288 -228 -5380
rect 48 -7086 78 8820
rect 266 4436 276 4488
rect 328 4436 338 4488
rect 23250 3636 23260 3654
rect 21442 3606 23260 3636
rect 23250 3602 23260 3606
rect 23312 3602 23322 3654
rect 695 -619 705 -567
rect 757 -619 767 -567
rect 23278 -4716 23288 -4714
rect 20592 -4760 23288 -4716
rect 23278 -4766 23288 -4760
rect 23340 -4766 23350 -4714
rect 242 -5394 252 -5342
rect 304 -5394 314 -5342
rect 120 -7058 130 -7006
rect 182 -7058 192 -7006
rect 48 -7116 138 -7086
rect 23530 -7098 23560 9410
rect 23610 -4764 23620 -4712
rect 23672 -4764 23682 -4712
rect 696 -14821 706 -14769
rect 758 -14821 768 -14769
rect 20604 -18966 23372 -18924
rect 23362 -18976 23372 -18966
rect 23424 -18976 23434 -18924
rect 232 -19598 242 -19546
rect 294 -19598 304 -19546
rect 120 -21258 130 -21206
rect 182 -21258 192 -21206
rect -258 -21318 146 -21288
rect 23620 -21290 23650 -4764
rect 23680 -18974 23690 -18922
rect 23742 -18974 23752 -18922
rect -258 -21320 -228 -21318
rect 23586 -21328 23650 -21290
rect 696 -29031 706 -28979
rect 758 -29031 768 -28979
rect 20600 -33208 23190 -33160
rect 23180 -33212 23190 -33208
rect 23242 -33212 23252 -33160
rect 238 -33802 248 -33750
rect 300 -33802 310 -33750
rect 120 -35466 130 -35414
rect 182 -35466 192 -35414
rect -678 -35528 140 -35496
rect 23690 -35500 23720 -18974
rect 23824 -33212 23834 -33160
rect 23886 -33212 23896 -33160
rect -678 -35532 -648 -35528
rect 23582 -35538 23720 -35500
rect 696 -43233 706 -43181
rect 758 -43233 768 -43181
rect 20580 -46908 24124 -46858
rect -126 -47932 -116 -47918
rect -142 -47974 -116 -47932
rect -60 -47932 -50 -47918
rect -60 -47974 278 -47932
rect -142 -47988 278 -47974
rect 120 -49668 130 -49616
rect 182 -49668 192 -49616
rect 23800 -49700 23810 -49688
rect -1090 -49730 134 -49700
rect 23588 -49740 23810 -49700
rect 23862 -49740 23872 -49688
rect 4572 -56558 4618 -56194
rect 24092 -56292 24124 -46908
rect 18244 -56358 24124 -56292
rect 3082 -56718 3092 -56654
rect 3156 -56718 3166 -56654
rect 2306 -57092 2316 -57004
rect 2302 -57120 2316 -57092
rect 2420 -57120 2430 -57004
rect 2302 -57650 2430 -57120
rect 4574 -57472 4616 -56558
rect 6018 -57366 6028 -57314
rect 6080 -57366 6090 -57314
rect 3826 -57520 4616 -57472
rect 3826 -57530 4614 -57520
rect 6030 -57556 6060 -57366
rect 18244 -57552 18274 -56358
rect 21694 -57110 21704 -57046
rect 21768 -57110 21778 -57046
rect 1592 -57748 2430 -57650
rect 1592 -57750 2426 -57748
rect 1592 -57906 1692 -57750
rect 3836 -58540 3846 -58476
rect 3910 -58540 3920 -58476
rect 3654 -59456 3730 -59444
rect 3650 -59522 3660 -59456
rect 3724 -59498 3734 -59456
rect 3842 -59490 3904 -59438
rect 3842 -59492 16664 -59490
rect 3724 -59522 3762 -59498
rect 3654 -59534 3762 -59522
rect 3720 -59864 3762 -59534
rect 3832 -59556 3842 -59492
rect 3906 -59554 16664 -59492
rect 3906 -59556 3916 -59554
rect 3842 -59938 3904 -59556
rect 5010 -59640 5044 -59554
rect 5322 -59642 5356 -59554
rect 5428 -59640 5462 -59554
rect 5742 -59642 5776 -59554
rect 5850 -59642 5884 -59554
rect 6158 -59642 6192 -59554
rect 6266 -59642 6300 -59554
rect 6578 -59642 6612 -59554
rect 6684 -59642 6718 -59554
rect 6994 -59642 7028 -59554
rect 7102 -59642 7136 -59554
rect 7412 -59642 7446 -59554
rect 7520 -59642 7554 -59554
rect 7832 -59642 7866 -59554
rect 7938 -59642 7972 -59554
rect 8250 -59642 8284 -59554
rect 8358 -59638 8392 -59554
rect 8664 -59642 8698 -59554
rect 8776 -59642 8810 -59554
rect 9084 -59642 9118 -59554
rect 9192 -59642 9226 -59554
rect 9502 -59642 9536 -59554
rect 9610 -59642 9644 -59554
rect 9922 -59642 9956 -59554
rect 10030 -59642 10064 -59554
rect 10340 -59642 10374 -59554
rect 10446 -59642 10480 -59554
rect 10758 -59642 10792 -59554
rect 10866 -59640 10900 -59554
rect 11176 -59642 11210 -59554
rect 11284 -59642 11318 -59554
rect 11594 -59642 11628 -59554
rect 11700 -59642 11734 -59554
rect 12010 -59642 12044 -59554
rect 12120 -59642 12154 -59554
rect 12430 -59642 12464 -59554
rect 12538 -59642 12572 -59554
rect 12846 -59644 12880 -59554
rect 12952 -59640 12986 -59554
rect 13264 -59642 13298 -59554
rect 13372 -59642 13406 -59554
rect 13682 -59642 13716 -59554
rect 13790 -59642 13824 -59554
rect 14098 -59642 14132 -59554
rect 14210 -59640 14244 -59554
rect 14518 -59642 14552 -59554
rect 14630 -59640 14664 -59554
rect 14938 -59642 14972 -59554
rect 15046 -59642 15080 -59554
rect 15354 -59640 15388 -59554
rect 15464 -59642 15498 -59554
rect 15774 -59642 15808 -59554
rect 15882 -59642 15916 -59554
rect 16192 -59642 16226 -59554
rect 16298 -59646 16332 -59554
rect 16608 -59650 16642 -59554
rect 5064 -59754 16600 -59718
rect 5138 -59996 5174 -59754
rect 6864 -59996 6900 -59754
rect 8964 -59996 9000 -59754
rect 11482 -59996 11518 -59754
rect 5094 -60030 13550 -59996
rect 5022 -60114 5062 -60072
rect 5332 -60080 5370 -60070
rect 5332 -60114 5372 -60080
rect 5442 -60086 5480 -60072
rect 5022 -60276 5056 -60114
rect 5146 -60176 5156 -60124
rect 5208 -60176 5218 -60124
rect 5338 -60276 5372 -60114
rect 5436 -60114 5480 -60086
rect 5436 -60276 5470 -60114
rect 5748 -60116 5792 -60066
rect 5856 -60080 5900 -60066
rect 5854 -60116 5900 -60080
rect 5572 -60172 5582 -60120
rect 5634 -60172 5644 -60120
rect 5754 -60276 5788 -60116
rect 5854 -60276 5888 -60116
rect 6168 -60118 6212 -60068
rect 6276 -60112 6320 -60062
rect 6002 -60172 6012 -60120
rect 6064 -60172 6074 -60120
rect 6170 -60276 6204 -60118
rect 6280 -60276 6314 -60112
rect 6588 -60114 6632 -60064
rect 6696 -60082 6740 -60060
rect 7010 -60062 7054 -60060
rect 6690 -60110 6740 -60082
rect 7004 -60110 7054 -60062
rect 6412 -60174 6422 -60122
rect 6474 -60174 6484 -60122
rect 6596 -60276 6630 -60114
rect 6690 -60276 6724 -60110
rect 7004 -60112 7048 -60110
rect 6836 -60178 6846 -60126
rect 6898 -60178 6908 -60126
rect 7004 -60276 7038 -60112
rect 7114 -60114 7158 -60064
rect 7422 -60114 7466 -60064
rect 7530 -60092 7574 -60064
rect 7842 -60084 7886 -60062
rect 7524 -60114 7574 -60092
rect 7838 -60112 7886 -60084
rect 7948 -60110 7992 -60060
rect 7114 -60276 7148 -60114
rect 7256 -60174 7266 -60122
rect 7318 -60174 7328 -60122
rect 7430 -60276 7464 -60114
rect 7524 -60276 7558 -60114
rect 7678 -60180 7688 -60128
rect 7740 -60180 7750 -60128
rect 7838 -60276 7872 -60112
rect 7948 -60276 7982 -60110
rect 8258 -60112 8302 -60062
rect 8366 -60096 8410 -60060
rect 8364 -60110 8410 -60096
rect 8678 -60098 8722 -60060
rect 8676 -60110 8722 -60098
rect 8784 -60110 8828 -60060
rect 9096 -60108 9140 -60060
rect 9506 -60068 9550 -60062
rect 9094 -60110 9140 -60108
rect 8086 -60168 8096 -60116
rect 8148 -60168 8158 -60116
rect 8260 -60276 8294 -60112
rect 8364 -60276 8398 -60110
rect 8512 -60170 8522 -60118
rect 8574 -60170 8584 -60118
rect 8676 -60276 8710 -60110
rect 8788 -60276 8822 -60110
rect 8926 -60176 8936 -60124
rect 8988 -60176 8998 -60124
rect 9094 -60276 9128 -60110
rect 9500 -60112 9550 -60068
rect 9814 -60110 9858 -60060
rect 9924 -60070 9968 -60062
rect 9500 -60252 9534 -60112
rect 9666 -60176 9676 -60124
rect 9728 -60176 9738 -60124
rect 9814 -60252 9848 -60110
rect 9918 -60112 9968 -60070
rect 10232 -60110 10276 -60060
rect 10342 -60110 10386 -60060
rect 9918 -60252 9952 -60112
rect 10066 -60168 10076 -60116
rect 10128 -60168 10138 -60116
rect 10236 -60252 10270 -60110
rect 10342 -60252 10376 -60110
rect 10652 -60112 10696 -60062
rect 10760 -60112 10804 -60062
rect 11068 -60074 11112 -60062
rect 11068 -60112 11116 -60074
rect 11176 -60080 11220 -60060
rect 11176 -60110 11222 -60080
rect 10476 -60174 10486 -60122
rect 10538 -60174 10548 -60122
rect 10652 -60252 10686 -60112
rect 10768 -60252 10802 -60112
rect 10900 -60174 10910 -60122
rect 10962 -60174 10972 -60122
rect 11082 -60252 11116 -60112
rect 11188 -60252 11222 -60110
rect 11486 -60112 11530 -60062
rect 11596 -60110 11640 -60060
rect 11904 -60070 11938 -60068
rect 11322 -60174 11332 -60122
rect 11384 -60174 11394 -60122
rect 11494 -60252 11528 -60112
rect 11598 -60250 11632 -60110
rect 11904 -60116 11942 -60070
rect 12012 -60110 12056 -60060
rect 12316 -60062 12350 -60058
rect 11732 -60176 11742 -60124
rect 11794 -60176 11804 -60124
rect 11598 -60252 11676 -60250
rect 11904 -60252 11938 -60116
rect 12020 -60252 12054 -60110
rect 12316 -60112 12368 -60062
rect 12430 -60110 12474 -60060
rect 12740 -60082 12784 -60062
rect 12150 -60172 12160 -60120
rect 12212 -60172 12222 -60120
rect 12316 -60252 12350 -60112
rect 12436 -60252 12470 -60110
rect 12740 -60112 12788 -60082
rect 12850 -60110 12894 -60060
rect 13160 -60062 13194 -60058
rect 13276 -60062 13310 -60060
rect 13586 -60062 13620 -60060
rect 12572 -60170 12582 -60118
rect 12634 -60170 12644 -60118
rect 12754 -60252 12788 -60112
rect 12854 -60252 12888 -60110
rect 13158 -60112 13202 -60062
rect 13266 -60112 13310 -60062
rect 13576 -60112 13620 -60062
rect 12992 -60178 13002 -60126
rect 13054 -60178 13064 -60126
rect 13160 -60252 13194 -60112
rect 13276 -60252 13310 -60112
rect 13410 -60174 13420 -60122
rect 13472 -60174 13482 -60122
rect 13586 -60250 13620 -60112
rect 21692 -60250 21702 -60228
rect 13586 -60252 21702 -60250
rect 5018 -60324 9154 -60276
rect 9500 -60292 21702 -60252
rect 21766 -60250 21776 -60228
rect 21766 -60292 21790 -60250
rect 9500 -60300 21790 -60292
rect 3064 -60366 3166 -60362
rect 3064 -60430 3084 -60366
rect 3148 -60390 3166 -60366
rect 5020 -60390 5064 -60324
rect 3148 -60430 5064 -60390
rect 3064 -60434 5064 -60430
rect 3064 -60438 3166 -60434
<< via1 >>
rect -258 -5380 -206 -5328
rect -676 -19582 -624 -19530
rect -1084 -33752 -1032 -33700
rect 276 4436 328 4488
rect 23260 3602 23312 3654
rect 705 -619 757 -567
rect 23288 -4766 23340 -4714
rect 252 -5394 304 -5342
rect 130 -7058 182 -7006
rect 23620 -4764 23672 -4712
rect 706 -14821 758 -14769
rect 23372 -18976 23424 -18924
rect 242 -19598 294 -19546
rect 130 -21258 182 -21206
rect 23690 -18974 23742 -18922
rect 706 -29031 758 -28979
rect 23190 -33212 23242 -33160
rect 248 -33802 300 -33750
rect 130 -35466 182 -35414
rect 23834 -33212 23886 -33160
rect 706 -43233 758 -43181
rect -116 -47974 -60 -47918
rect 130 -49668 182 -49616
rect 23810 -49740 23862 -49688
rect 3092 -56718 3156 -56654
rect 2316 -57120 2420 -57004
rect 6028 -57366 6080 -57314
rect 21704 -57110 21768 -57046
rect 3846 -58540 3910 -58476
rect 3660 -59522 3724 -59456
rect 3842 -59556 3906 -59492
rect 5156 -60176 5208 -60124
rect 5582 -60172 5634 -60120
rect 6012 -60172 6064 -60120
rect 6422 -60174 6474 -60122
rect 6846 -60178 6898 -60126
rect 7266 -60174 7318 -60122
rect 7688 -60180 7740 -60128
rect 8096 -60168 8148 -60116
rect 8522 -60170 8574 -60118
rect 8936 -60176 8988 -60124
rect 9676 -60176 9728 -60124
rect 10076 -60168 10128 -60116
rect 10486 -60174 10538 -60122
rect 10910 -60174 10962 -60122
rect 11332 -60174 11384 -60122
rect 11742 -60176 11794 -60124
rect 12160 -60172 12212 -60120
rect 12582 -60170 12634 -60118
rect 13002 -60178 13054 -60126
rect 13420 -60174 13472 -60122
rect 21702 -60292 21766 -60228
rect 3084 -60430 3148 -60366
<< metal2 >>
rect 276 4488 328 4498
rect -2732 4466 276 4484
rect -2734 4436 276 4466
rect -2734 4434 328 4436
rect -2734 -60168 -2686 4434
rect 276 4426 328 4434
rect 748 -557 788 803
rect 705 -567 788 -557
rect 757 -619 788 -567
rect 705 -623 788 -619
rect 705 -629 757 -623
rect -258 -5328 -206 -5318
rect 252 -5342 304 -5332
rect -206 -5380 252 -5346
rect -258 -5390 -206 -5380
rect 252 -5404 304 -5394
rect -1260 -7002 -1204 -6992
rect 130 -7004 182 -6996
rect -1204 -7006 182 -7004
rect -1204 -7058 130 -7006
rect -1260 -7068 -1204 -7058
rect 130 -7068 182 -7058
rect 750 -14759 790 -13394
rect 706 -14769 790 -14759
rect 758 -14820 790 -14769
rect 706 -14831 758 -14821
rect -676 -19530 -624 -19520
rect 242 -19546 294 -19536
rect -624 -19580 242 -19550
rect -676 -19592 -624 -19582
rect 242 -19608 294 -19598
rect -1272 -21204 -1216 -21194
rect -1276 -21260 -1272 -21208
rect 130 -21206 182 -21196
rect -1216 -21258 130 -21208
rect -1216 -21260 182 -21258
rect -1276 -21262 182 -21260
rect -1272 -21270 -1216 -21262
rect 130 -21268 182 -21262
rect 750 -28969 790 -27603
rect 706 -28979 790 -28969
rect 758 -29029 790 -28979
rect 706 -29041 758 -29031
rect -1084 -33700 -1032 -33690
rect 248 -33750 300 -33740
rect -1032 -33752 248 -33750
rect -1084 -33762 248 -33752
rect -1074 -33794 248 -33762
rect 248 -33812 300 -33802
rect -1288 -35412 -1232 -35402
rect 130 -35414 182 -35404
rect -1232 -35466 130 -35416
rect -1232 -35468 182 -35466
rect -1288 -35470 182 -35468
rect -1288 -35478 -1232 -35470
rect 130 -35476 182 -35470
rect 750 -43171 790 -41812
rect 706 -43181 790 -43171
rect 758 -43233 790 -43181
rect 706 -43238 790 -43233
rect 706 -43243 758 -43238
rect -116 -47918 -60 -47908
rect -116 -47984 -60 -47974
rect -1266 -49614 -1210 -49604
rect -1268 -49670 -1266 -49620
rect 130 -49616 182 -49606
rect -1210 -49668 130 -49620
rect -1210 -49670 182 -49668
rect -1268 -49674 182 -49670
rect -1266 -49680 -1210 -49674
rect 130 -49678 182 -49674
rect -116 -49948 -60 -49938
rect -116 -50014 -60 -50004
rect -114 -57310 -62 -50014
rect 2289 -55554 2441 13391
rect 22589 -51048 23031 8837
rect 23260 3654 23312 3664
rect 23312 3606 24956 3642
rect 23260 3592 23312 3602
rect 23288 -4714 23340 -4704
rect 23620 -4712 23672 -4702
rect 23340 -4762 23620 -4714
rect 23288 -4776 23340 -4766
rect 23620 -4774 23672 -4764
rect 23372 -18924 23424 -18914
rect 23690 -18922 23742 -18912
rect 23424 -18974 23690 -18926
rect 23424 -18976 23742 -18974
rect 23372 -18986 23424 -18976
rect 23690 -18984 23742 -18976
rect 23190 -33160 23242 -33150
rect 23834 -33160 23886 -33150
rect 23242 -33212 23834 -33160
rect 23190 -33222 23242 -33212
rect 23832 -33222 23886 -33212
rect 23832 -49678 23862 -33222
rect 23810 -49688 23862 -49678
rect 23810 -49750 23862 -49740
rect 2289 -55599 2442 -55554
rect 2290 -57004 2442 -55599
rect 3092 -56654 3156 -56644
rect 3092 -56728 3156 -56718
rect 2290 -57120 2316 -57004
rect 2420 -57120 2442 -57004
rect 21704 -57046 21768 -57036
rect 21704 -57120 21768 -57110
rect 2290 -57146 2442 -57120
rect 6028 -57310 6080 -57304
rect -114 -57314 6084 -57310
rect -114 -57366 6028 -57314
rect 6080 -57366 6084 -57314
rect 6028 -57376 6080 -57366
rect 3846 -58476 3910 -58466
rect 3846 -58550 3910 -58540
rect 3660 -59456 3724 -59446
rect 3660 -59532 3724 -59522
rect 3842 -59492 3906 -59482
rect 3842 -59566 3906 -59556
rect 5156 -60124 5208 -60114
rect -2734 -60176 5156 -60168
rect 5582 -60120 5634 -60110
rect 5208 -60172 5582 -60168
rect 6012 -60120 6064 -60110
rect 5634 -60172 6012 -60168
rect 6422 -60122 6474 -60112
rect 6064 -60172 6422 -60168
rect 5208 -60174 6422 -60172
rect 6846 -60126 6898 -60116
rect 6474 -60174 6846 -60168
rect 5208 -60176 6846 -60174
rect -2734 -60178 6846 -60176
rect 7266 -60122 7318 -60112
rect 8096 -60116 8148 -60106
rect 6898 -60174 7266 -60168
rect 7688 -60128 7740 -60118
rect 7318 -60174 7688 -60168
rect 6898 -60178 7688 -60174
rect -2734 -60180 7688 -60178
rect 8522 -60118 8574 -60108
rect 7740 -60170 8522 -60168
rect 8936 -60124 8988 -60114
rect 8574 -60170 8936 -60168
rect 7740 -60176 8936 -60170
rect 9676 -60124 9728 -60114
rect 8988 -60176 8998 -60168
rect 7740 -60180 8998 -60176
rect -2734 -60214 8998 -60180
rect 9666 -60176 9676 -60168
rect 10076 -60116 10128 -60106
rect 10486 -60122 10538 -60112
rect 9728 -60174 10486 -60168
rect 10910 -60122 10962 -60112
rect 10538 -60174 10910 -60168
rect 11332 -60122 11384 -60112
rect 10962 -60174 11332 -60168
rect 11742 -60124 11794 -60114
rect 11384 -60174 11742 -60168
rect 9728 -60176 11742 -60174
rect 12160 -60120 12212 -60110
rect 11794 -60172 12160 -60168
rect 12582 -60118 12634 -60108
rect 12212 -60170 12582 -60168
rect 13002 -60126 13054 -60116
rect 12634 -60170 13002 -60168
rect 12212 -60172 13002 -60170
rect 11794 -60176 13002 -60172
rect 9666 -60178 13002 -60176
rect 13420 -60122 13472 -60112
rect 13054 -60174 13420 -60168
rect 24896 -60132 24954 3606
rect 16098 -60164 24954 -60132
rect 16098 -60168 24950 -60164
rect 13472 -60174 24950 -60168
rect 13054 -60178 24950 -60174
rect 9666 -60180 24950 -60178
rect 9666 -60214 16176 -60180
rect 21702 -60228 21766 -60218
rect 21702 -60302 21766 -60292
rect 3084 -60366 3148 -60356
rect 3084 -60440 3148 -60430
<< via2 >>
rect -1260 -7058 -1204 -7002
rect -1272 -21260 -1216 -21204
rect -1288 -35468 -1232 -35412
rect -116 -47974 -60 -47918
rect -1266 -49670 -1210 -49614
rect -116 -50004 -60 -49948
rect 3092 -56718 3156 -56654
rect 21704 -57110 21768 -57046
rect 3846 -58540 3910 -58476
rect 3660 -59522 3724 -59456
rect 3842 -59556 3906 -59492
rect 21702 -60292 21766 -60228
rect 3084 -60430 3148 -60366
<< metal3 >>
rect -1270 -7002 -1194 -6997
rect -1270 -7008 -1260 -7002
rect -1276 -7058 -1260 -7008
rect -1204 -7058 -1194 -7002
rect -1276 -21199 -1194 -7058
rect -1282 -21204 -1194 -21199
rect -1282 -21260 -1272 -21204
rect -1216 -21260 -1194 -21204
rect -1282 -21265 -1194 -21260
rect -1276 -35407 -1194 -21265
rect -1298 -35412 -1194 -35407
rect -1298 -35468 -1288 -35412
rect -1232 -35468 -1194 -35412
rect -1298 -35473 -1194 -35468
rect -1276 -49614 -1194 -35473
rect -126 -47916 -50 -47913
rect -1276 -49670 -1266 -49614
rect -1210 -49670 -1194 -49614
rect -150 -47918 -50 -47916
rect -150 -47974 -116 -47918
rect -60 -47974 -50 -47918
rect -150 -47979 -50 -47974
rect -1276 -49675 -1200 -49670
rect -150 -49943 -52 -47979
rect -150 -49948 -50 -49943
rect -150 -50004 -116 -49948
rect -60 -50004 -50 -49948
rect -150 -50009 -50 -50004
rect -150 -50010 -52 -50009
rect 335 -56390 490 14085
rect 1238 13450 1348 13486
rect 334 -56504 490 -56390
rect 334 -58970 530 -56504
rect 3074 -56654 3224 -56602
rect 3074 -56718 3092 -56654
rect 3156 -56718 3224 -56654
rect 3074 -56724 3224 -56718
rect 21682 -57046 21810 -56996
rect 21682 -57110 21704 -57046
rect 21768 -57110 21810 -57046
rect 21682 -57126 21810 -57110
rect 3820 -58476 3920 -58448
rect 3820 -58540 3846 -58476
rect 3910 -58540 3920 -58476
rect 3820 -58548 3920 -58540
rect 3250 -59272 3538 -58964
rect 3250 -59418 3732 -59272
rect 3250 -59456 3734 -59418
rect 3250 -59480 3660 -59456
rect 3250 -60056 3538 -59480
rect 3650 -59522 3660 -59480
rect 3724 -59522 3734 -59456
rect 3650 -59527 3734 -59522
rect 3822 -59492 3922 -59422
rect 3822 -59556 3842 -59492
rect 3906 -59556 3922 -59492
rect 3822 -59560 3922 -59556
rect 3832 -59561 3916 -59560
rect 21680 -60228 21782 -60210
rect 21680 -60292 21702 -60228
rect 21766 -60292 21782 -60228
rect 21680 -60308 21782 -60292
rect 3052 -60366 3178 -60336
rect 3052 -60430 3084 -60366
rect 3148 -60430 3178 -60366
rect 3052 -60442 3178 -60430
<< via3 >>
rect 3092 -56718 3156 -56654
rect 21704 -57110 21768 -57046
rect 3846 -58540 3910 -58476
rect 3842 -59556 3906 -59492
rect 21702 -60292 21766 -60228
rect 3084 -60430 3148 -60366
<< metal4 >>
rect 1279 -52251 1350 13486
rect 3086 -56654 3158 -56648
rect 3086 -56718 3092 -56654
rect 3156 -56718 3158 -56654
rect 3086 -60130 3158 -56718
rect 21700 -57045 21768 -57042
rect 21700 -57046 21769 -57045
rect 21700 -57110 21704 -57046
rect 21768 -57110 21769 -57046
rect 21700 -57111 21769 -57110
rect 3845 -58476 3911 -58475
rect 3842 -58540 3846 -58476
rect 3910 -58540 3911 -58476
rect 3842 -58541 3911 -58540
rect 3842 -59491 3902 -58541
rect 3841 -59492 3907 -59491
rect 3841 -59556 3842 -59492
rect 3906 -59556 3907 -59492
rect 3841 -59557 3907 -59556
rect 3084 -60365 3158 -60130
rect 21700 -60228 21768 -57111
rect 21700 -60292 21702 -60228
rect 21766 -60292 21768 -60228
rect 21700 -60296 21768 -60292
rect 3083 -60366 3158 -60365
rect 3083 -60430 3084 -60366
rect 3148 -60430 3158 -60366
rect 3083 -60431 3149 -60430
use fb  fb_0
timestamp 1662983156
transform 1 0 -45844 0 1 -51192
box 46324 -8198 69992 -5432
use sky130_fd_pr__nfet_01v8_lvt_8PSHEW  sky130_fd_pr__nfet_01v8_lvt_8PSHEW_0
timestamp 1662988209
transform 1 0 3819 0 1 -59732
box -211 -338 211 338
use sky130_fd_pr__nfet_01v8_lvt_72NHPP  sky130_fd_pr__nfet_01v8_lvt_72NHPP_0
timestamp 1662988209
transform 0 1 7077 -1 0 -60093
box -211 -2191 211 2191
use sky130_fd_pr__nfet_01v8_lvt_72NHPP  sky130_fd_pr__nfet_01v8_lvt_72NHPP_1
timestamp 1662988209
transform 0 1 11559 -1 0 -60093
box -211 -2191 211 2191
use sky130_fd_pr__nfet_01v8_lvt_XA5MKQ  sky130_fd_pr__nfet_01v8_lvt_XA5MKQ_0
timestamp 1662988209
transform 0 1 10827 -1 0 -59659
box -211 -5953 211 5953
use stage0  stage0_0
timestamp 1662974608
transform 1 0 18 0 1 5376
box 0 -5324 26310 8797
use stage1  stage1_0
timestamp 1662978535
transform 1 0 20 0 1 -8826
box 0 -5324 26310 8797
use stage1  stage1_1
timestamp 1662978535
transform 1 0 20 0 1 -23028
box 0 -5324 26310 8797
use stage1  stage1_2
timestamp 1662978535
transform 1 0 20 0 1 -37238
box 0 -5324 26310 8797
use stage1  stage1_3
timestamp 1662978535
transform 1 0 20 0 1 -51440
box 0 -5324 26310 8797
<< labels >>
rlabel space 2274 8444 2441 13391 0 vdd
rlabel space 304 8136 490 14085 0 vss
rlabel space 968 13660 1017 14026 0 Iref
rlabel metal3 1238 13450 1348 13486 0 vref
rlabel metal2 -1204 -7058 130 -7004 0 vc
rlabel metal2 -114 -57366 -62 -50004 0 vout5p
rlabel space 18244 -58136 18274 -56292 0 vout5n
rlabel space 128 7086 4168 7116 0 vinp
rlabel space 128 7026 4078 7056 0 vinn
rlabel metal1 13586 -60300 21702 -60250 0 vin0n
rlabel metal1 5020 -60434 5064 -60276 0 vin0p
<< end >>
