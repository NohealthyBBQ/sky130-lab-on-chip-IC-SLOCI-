magic
tech sky130A
magscale 1 2
timestamp 1662405622
<< pwell >>
rect 7710 2035 7715 2140
<< locali >>
rect 6405 3125 6675 3160
rect 7100 3125 7370 3160
rect 7840 3125 8110 3160
rect 6410 1935 6680 1970
rect 7135 1935 7405 1970
rect 7840 1935 8110 1970
rect 6410 1750 6680 1785
rect 7145 1750 7415 1785
rect 7830 1750 8100 1785
rect 6405 1435 6675 1470
rect 7145 1435 7415 1470
rect 7850 1435 8120 1470
<< metal1 >>
rect 5155 8490 6315 8510
rect 5155 8095 5175 8490
rect 6295 8095 6315 8490
rect 5155 8075 6315 8095
rect 8200 8490 9360 8510
rect 8200 8095 8220 8490
rect 9340 8095 9360 8490
rect 8200 8075 9360 8095
rect 5000 3125 9520 3185
rect 6720 2085 6780 3125
rect 6810 3050 6895 3060
rect 6810 2995 6820 3050
rect 6885 3000 7010 3050
rect 6885 2995 6895 3000
rect 6810 2990 6895 2995
rect 6930 2965 7010 2970
rect 6930 2956 6940 2965
rect 6810 2910 6940 2956
rect 7000 2910 7010 2965
rect 6810 2905 7010 2910
rect 6930 2900 7010 2905
rect 6810 2865 6895 2875
rect 6810 2810 6820 2865
rect 6885 2860 6895 2865
rect 6885 2810 7010 2860
rect 6810 2805 6895 2810
rect 6930 2770 7010 2780
rect 6930 2762 6940 2770
rect 6810 2715 6940 2762
rect 7000 2715 7010 2770
rect 6810 2710 7010 2715
rect 6930 2705 7010 2710
rect 6810 2670 6895 2680
rect 6810 2615 6820 2670
rect 6885 2620 7010 2670
rect 6885 2615 6895 2620
rect 6810 2605 6895 2615
rect 6930 2580 7010 2590
rect 6930 2571 6940 2580
rect 6810 2525 6940 2571
rect 7000 2525 7010 2580
rect 6810 2520 7010 2525
rect 6930 2515 7010 2520
rect 6810 2480 6895 2490
rect 6810 2425 6820 2480
rect 6885 2475 6895 2480
rect 6885 2425 7010 2475
rect 6810 2415 6895 2425
rect 6930 2385 7010 2395
rect 6930 2378 6940 2385
rect 6810 2330 6940 2378
rect 7000 2330 7010 2385
rect 6810 2325 7010 2330
rect 6930 2320 7010 2325
rect 6810 2285 6895 2295
rect 6810 2230 6820 2285
rect 6885 2235 7010 2285
rect 6885 2230 6895 2235
rect 6810 2220 6895 2230
rect 6930 2195 7010 2205
rect 6930 2186 6940 2195
rect 6810 2140 6940 2186
rect 7000 2140 7010 2195
rect 7040 2175 7100 3125
rect 7420 2175 7480 3125
rect 7625 3050 7710 3060
rect 7510 3000 7635 3050
rect 7625 2995 7635 3000
rect 7700 2995 7710 3050
rect 7625 2990 7710 2995
rect 7510 2965 7590 2970
rect 7510 2910 7520 2965
rect 7580 2956 7590 2965
rect 7580 2910 7710 2956
rect 7510 2905 7710 2910
rect 7510 2900 7590 2905
rect 7625 2865 7710 2875
rect 7625 2860 7635 2865
rect 7510 2810 7635 2860
rect 7700 2810 7710 2865
rect 7625 2805 7710 2810
rect 7510 2770 7590 2780
rect 7510 2715 7520 2770
rect 7580 2761 7590 2770
rect 7580 2715 7710 2761
rect 7510 2710 7710 2715
rect 7510 2705 7590 2710
rect 7625 2670 7710 2680
rect 7510 2620 7635 2670
rect 7625 2615 7635 2620
rect 7700 2615 7710 2670
rect 7625 2605 7710 2615
rect 7510 2580 7590 2590
rect 7510 2525 7520 2580
rect 7580 2571 7590 2580
rect 7580 2525 7710 2571
rect 7510 2520 7710 2525
rect 7510 2515 7590 2520
rect 7625 2480 7710 2490
rect 7625 2475 7635 2480
rect 7510 2425 7635 2475
rect 7700 2425 7710 2480
rect 7625 2415 7710 2425
rect 7510 2385 7590 2390
rect 7510 2330 7520 2385
rect 7580 2376 7590 2385
rect 7580 2330 7710 2376
rect 7510 2325 7710 2330
rect 7510 2320 7590 2325
rect 7625 2285 7710 2295
rect 7510 2235 7635 2285
rect 7625 2230 7635 2235
rect 7700 2230 7710 2285
rect 7625 2220 7710 2230
rect 7510 2195 7590 2205
rect 6810 2135 7010 2140
rect 6930 2130 7010 2135
rect 7510 2140 7520 2195
rect 7580 2185 7590 2195
rect 7580 2140 7710 2185
rect 7510 2135 7710 2140
rect 7510 2130 7590 2135
rect 6810 2095 6895 2105
rect 6810 2040 6820 2095
rect 6885 2090 6895 2095
rect 7625 2095 7710 2105
rect 7625 2090 7635 2095
rect 6885 2040 7015 2090
rect 7505 2040 7635 2090
rect 7700 2040 7710 2095
rect 7740 2085 7800 3125
rect 6810 2035 6895 2040
rect 7625 2035 7710 2040
rect 5165 1980 6315 2000
rect 5165 1585 5185 1980
rect 6295 1585 6315 1980
rect 8205 1980 9350 1995
rect 6810 1715 7010 1725
rect 5165 1565 6315 1585
rect 6730 1450 6780 1645
rect 6810 1640 6820 1715
rect 7000 1640 7010 1715
rect 7510 1715 7710 1725
rect 6810 1630 7010 1640
rect 6810 1580 7010 1590
rect 6810 1515 6820 1580
rect 7000 1515 7010 1580
rect 6810 1505 7010 1515
rect 7040 1450 7090 1645
rect 6730 1400 7090 1450
rect 7430 1450 7480 1645
rect 7510 1640 7520 1715
rect 7700 1640 7710 1715
rect 7510 1630 7710 1640
rect 7510 1580 7710 1590
rect 7510 1515 7520 1580
rect 7700 1515 7710 1580
rect 7510 1505 7710 1515
rect 7740 1450 7790 1645
rect 8205 1585 8225 1980
rect 9335 1585 9350 1980
rect 8205 1565 9350 1585
rect 7430 1400 7790 1450
<< via1 >>
rect 5175 8095 6295 8490
rect 8220 8095 9340 8490
rect 6820 2995 6885 3050
rect 6940 2910 7000 2965
rect 6820 2810 6885 2865
rect 6940 2715 7000 2770
rect 6820 2615 6885 2670
rect 6940 2525 7000 2580
rect 6820 2425 6885 2480
rect 6940 2330 7000 2385
rect 6820 2230 6885 2285
rect 6940 2140 7000 2195
rect 7635 2995 7700 3050
rect 7520 2910 7580 2965
rect 7635 2810 7700 2865
rect 7520 2715 7580 2770
rect 7635 2615 7700 2670
rect 7520 2525 7580 2580
rect 7635 2425 7700 2480
rect 7520 2330 7580 2385
rect 7635 2230 7700 2285
rect 7520 2140 7580 2195
rect 6820 2040 6885 2095
rect 7635 2040 7700 2095
rect 5185 1585 6295 1980
rect 6820 1640 7000 1715
rect 6820 1515 7000 1580
rect 7520 1640 7700 1715
rect 7520 1515 7700 1580
rect 8225 1585 9335 1980
<< metal2 >>
rect 5000 8490 9520 8510
rect 5000 8095 5175 8490
rect 6295 8095 8220 8490
rect 9340 8095 9520 8490
rect 5000 8070 9520 8095
rect 5000 3225 9520 3625
rect 6495 3050 6895 3225
rect 6495 2995 6820 3050
rect 6885 2995 6895 3050
rect 6495 2865 6895 2995
rect 7040 2975 7480 3065
rect 7625 3050 8025 3225
rect 7625 2995 7635 3050
rect 7700 2995 8025 3050
rect 6930 2965 7590 2975
rect 6930 2910 6940 2965
rect 7000 2910 7520 2965
rect 7580 2910 7590 2965
rect 6930 2900 7590 2910
rect 6495 2810 6820 2865
rect 6885 2810 6895 2865
rect 6495 2670 6895 2810
rect 7040 2780 7480 2900
rect 7625 2865 8025 2995
rect 7625 2810 7635 2865
rect 7700 2810 8025 2865
rect 6930 2770 7590 2780
rect 6930 2715 6940 2770
rect 7000 2715 7520 2770
rect 7580 2715 7590 2770
rect 6930 2705 7590 2715
rect 6495 2615 6820 2670
rect 6885 2615 6895 2670
rect 6495 2480 6895 2615
rect 7040 2590 7480 2705
rect 7625 2670 8025 2810
rect 7625 2615 7635 2670
rect 7700 2615 8025 2670
rect 6930 2580 7590 2590
rect 6930 2525 6940 2580
rect 7000 2525 7520 2580
rect 7580 2525 7590 2580
rect 6930 2515 7590 2525
rect 6495 2425 6820 2480
rect 6885 2425 6895 2480
rect 6495 2285 6895 2425
rect 7040 2395 7480 2515
rect 7625 2480 8025 2615
rect 7625 2425 7635 2480
rect 7700 2425 8025 2480
rect 6930 2385 7590 2395
rect 6930 2330 6940 2385
rect 7000 2330 7520 2385
rect 7580 2330 7590 2385
rect 6930 2320 7590 2330
rect 6495 2230 6820 2285
rect 6885 2230 6895 2285
rect 6495 2095 6895 2230
rect 7040 2205 7480 2320
rect 7625 2285 8025 2425
rect 7625 2230 7635 2285
rect 7700 2230 8025 2285
rect 6930 2195 7590 2205
rect 6930 2140 6940 2195
rect 7000 2140 7520 2195
rect 7580 2140 7590 2195
rect 6930 2130 7590 2140
rect 6495 2040 6820 2095
rect 6885 2040 6895 2095
rect 6495 2035 6895 2040
rect 5165 1980 6315 2000
rect 5165 1585 5185 1980
rect 6295 1585 6315 1980
rect 7040 1870 7480 2130
rect 7625 2095 8025 2230
rect 7625 2040 7635 2095
rect 7700 2040 8025 2095
rect 7625 2035 8025 2040
rect 8205 1980 9350 2000
rect 6715 1720 7805 1870
rect 6715 1715 7105 1720
rect 6715 1685 6820 1715
rect 6810 1640 6820 1685
rect 7000 1685 7105 1715
rect 7415 1715 7805 1720
rect 7415 1685 7520 1715
rect 7000 1640 7010 1685
rect 6810 1630 7010 1640
rect 7510 1640 7520 1685
rect 7700 1685 7805 1715
rect 7700 1640 7710 1685
rect 7510 1630 7710 1640
rect 5165 1565 6315 1585
rect 6810 1580 7010 1590
rect 6810 1515 6820 1580
rect 7000 1515 7010 1580
rect 6810 1505 7010 1515
rect 7510 1580 7710 1590
rect 7510 1515 7520 1580
rect 7700 1515 7710 1580
rect 8205 1585 8225 1980
rect 9335 1585 9350 1980
rect 8205 1570 9350 1585
rect 7510 1505 7710 1515
<< via2 >>
rect 5185 1585 6295 1980
rect 6820 1515 7000 1580
rect 7520 1515 7700 1580
rect 8225 1585 9335 1980
<< metal3 >>
rect 5165 1980 6315 2000
rect 5165 1585 5185 1980
rect 6295 1590 6315 1980
rect 8205 1980 9350 1995
rect 8205 1590 8225 1980
rect 6295 1585 7010 1590
rect 5165 1580 7010 1585
rect 5165 1515 6820 1580
rect 7000 1515 7010 1580
rect 5165 1410 7010 1515
rect 7510 1585 8225 1590
rect 9335 1585 9350 1980
rect 7510 1580 9350 1585
rect 7510 1515 7520 1580
rect 7700 1515 9350 1580
rect 7510 1410 9350 1515
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM1
timestamp 1662404926
transform 0 -1 6910 -1 0 2547
box -647 -310 647 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM2
timestamp 1662404926
transform 0 1 6910 -1 0 1611
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM3
timestamp 1662404926
transform 0 1 7610 -1 0 1611
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM4
timestamp 1662404926
transform 0 1 7610 -1 0 2547
box -647 -310 647 310
use sky130_fd_pr__res_high_po_5p73_YZEQ6M  XR1
timestamp 1662404926
transform 1 0 5739 0 1 5038
box -739 -3638 739 3638
use sky130_fd_pr__res_high_po_5p73_YZEQ6M  XR2
timestamp 1662404926
transform 1 0 8779 0 1 5038
box -739 -3638 739 3638
<< labels >>
rlabel metal1 7430 1400 7790 1450 1 INA
rlabel metal1 6730 1400 7090 1450 1 INB
rlabel metal1 5000 3125 9520 3185 1 BIAS
rlabel metal2 5000 3225 9520 3625 1 GND
rlabel metal2 6295 8075 8220 8510 1 VDD
rlabel metal3 5165 1410 6820 1585 1 OUTB
rlabel metal3 7700 1410 9350 1585 1 OUTA
rlabel locali 7145 1435 7415 1470 1 SUB
<< end >>
