magic
tech sky130A
magscale 1 2
timestamp 1662079606
use sky130_fd_pr__cap_mim_m3_1_EN3Q86  XC1
timestamp 1661639644
transform 1 0 -5538 0 1 2000
box -1750 -2240 1749 2240
use XM_actload2  XM_actload2_0
timestamp 1661870098
transform 1 0 5911 0 1 -2151
box -53 -53 2571 3173
use XM_cs  XM_cs_0
timestamp 1661891635
transform 1 0 8792 0 1 -2181
box -64 -53 2482 5609
use sky130_fd_pr__nfet_01v8_lvt_BRDQL2  XM_diff_n
timestamp 1661639644
transform 1 0 3416 0 1 13643
box -296 -2337 296 2337
use sky130_fd_pr__nfet_01v8_lvt_BRDQL2  XM_diff_n1
timestamp 1661639644
transform 1 0 5202 0 1 11615
box -296 -2337 296 2337
use XM_ppair  XM_ppair_0
timestamp 1662067076
transform 1 0 5958 0 1 8016
box -220 -1160 4440 828
use sky130_fd_pr__nfet_01v8_lvt_62X5LT  XM_tail
timestamp 1661892224
transform 1 0 3688 0 1 -89
box -1312 -657 1312 657
<< end >>
