magic
tech sky130A
magscale 1 2
timestamp 1662487295
<< error_p >>
rect -194 454 194 672
rect -194 18 194 236
rect -194 -418 194 -200
<< nwell >>
rect -194 454 194 854
rect -194 18 194 418
rect -194 -418 194 -18
rect -194 -854 194 -454
<< pmoslvt >>
rect -100 554 100 754
rect -100 118 100 318
rect -100 -318 100 -118
rect -100 -754 100 -554
<< pdiff >>
rect -158 742 -100 754
rect -158 566 -146 742
rect -112 566 -100 742
rect -158 554 -100 566
rect 100 742 158 754
rect 100 566 112 742
rect 146 566 158 742
rect 100 554 158 566
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -306 -146 -130
rect -112 -306 -100 -130
rect -158 -318 -100 -306
rect 100 -130 158 -118
rect 100 -306 112 -130
rect 146 -306 158 -130
rect 100 -318 158 -306
rect -158 -566 -100 -554
rect -158 -742 -146 -566
rect -112 -742 -100 -566
rect -158 -754 -100 -742
rect 100 -566 158 -554
rect 100 -742 112 -566
rect 146 -742 158 -566
rect 100 -754 158 -742
<< pdiffc >>
rect -146 566 -112 742
rect 112 566 146 742
rect -146 130 -112 306
rect 112 130 146 306
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -146 -742 -112 -566
rect 112 -742 146 -566
<< poly >>
rect -100 835 100 851
rect -100 801 -84 835
rect 84 801 100 835
rect -100 754 100 801
rect -100 507 100 554
rect -100 473 -84 507
rect 84 473 100 507
rect -100 457 100 473
rect -100 399 100 415
rect -100 365 -84 399
rect 84 365 100 399
rect -100 318 100 365
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -365 100 -318
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -415 100 -399
rect -100 -473 100 -457
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -100 -554 100 -507
rect -100 -801 100 -754
rect -100 -835 -84 -801
rect 84 -835 100 -801
rect -100 -851 100 -835
<< polycont >>
rect -84 801 84 835
rect -84 473 84 507
rect -84 365 84 399
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -84 -835 84 -801
<< locali >>
rect -100 801 -84 835
rect 84 801 100 835
rect -146 742 -112 758
rect -146 550 -112 566
rect 112 742 146 758
rect 112 550 146 566
rect -100 473 -84 507
rect 84 473 100 507
rect -100 365 -84 399
rect 84 365 100 399
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -322 -112 -306
rect 112 -130 146 -114
rect 112 -322 146 -306
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -507 -84 -473
rect 84 -507 100 -473
rect -146 -566 -112 -550
rect -146 -758 -112 -742
rect 112 -566 146 -550
rect 112 -758 146 -742
rect -100 -835 -84 -801
rect 84 -835 100 -801
<< viali >>
rect -84 801 84 835
rect -146 566 -112 742
rect 112 566 146 742
rect -84 473 84 507
rect -84 365 84 399
rect -146 130 -112 306
rect 112 130 146 306
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect -84 -399 84 -365
rect -84 -507 84 -473
rect -146 -742 -112 -566
rect 112 -742 146 -566
rect -84 -835 84 -801
<< metal1 >>
rect -96 835 96 841
rect -96 801 -84 835
rect 84 801 96 835
rect -96 795 96 801
rect -152 742 -106 754
rect -152 566 -146 742
rect -112 566 -106 742
rect -152 554 -106 566
rect 106 742 152 754
rect 106 566 112 742
rect 146 566 152 742
rect 106 554 152 566
rect -96 507 96 513
rect -96 473 -84 507
rect 84 473 96 507
rect -96 467 96 473
rect -96 399 96 405
rect -96 365 -84 399
rect 84 365 96 399
rect -96 359 96 365
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -306 -146 -130
rect -112 -306 -106 -130
rect -152 -318 -106 -306
rect 106 -130 152 -118
rect 106 -306 112 -130
rect 146 -306 152 -130
rect 106 -318 152 -306
rect -96 -365 96 -359
rect -96 -399 -84 -365
rect 84 -399 96 -365
rect -96 -405 96 -399
rect -96 -473 96 -467
rect -96 -507 -84 -473
rect 84 -507 96 -473
rect -96 -513 96 -507
rect -152 -566 -106 -554
rect -152 -742 -146 -566
rect -112 -742 -106 -566
rect -152 -754 -106 -742
rect 106 -566 152 -554
rect 106 -742 112 -566
rect 146 -742 152 -566
rect 106 -754 152 -742
rect -96 -801 96 -795
rect -96 -835 -84 -801
rect 84 -835 96 -801
rect -96 -841 96 -835
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 4 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
