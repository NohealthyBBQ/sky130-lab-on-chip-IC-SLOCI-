magic
tech sky130A
magscale 1 2
timestamp 1662726146
use sky130_fd_pr__nfet_01v8_lvt_4RBFJG  sky130_fd_pr__nfet_01v8_lvt_4RBFJG_0
timestamp 1662726146
transform 1 0 643 0 1 526
box -696 -579 696 579
<< end >>
