magic
tech sky130A
magscale 1 2
timestamp 1662486269
<< pwell >>
rect -1312 -1737 1312 1737
<< nmoslvt >>
rect -1116 927 -716 1527
rect -658 927 -258 1527
rect -200 927 200 1527
rect 258 927 658 1527
rect 716 927 1116 1527
rect -1116 109 -716 709
rect -658 109 -258 709
rect -200 109 200 709
rect 258 109 658 709
rect 716 109 1116 709
rect -1116 -709 -716 -109
rect -658 -709 -258 -109
rect -200 -709 200 -109
rect 258 -709 658 -109
rect 716 -709 1116 -109
rect -1116 -1527 -716 -927
rect -658 -1527 -258 -927
rect -200 -1527 200 -927
rect 258 -1527 658 -927
rect 716 -1527 1116 -927
<< ndiff >>
rect -1174 1515 -1116 1527
rect -1174 939 -1162 1515
rect -1128 939 -1116 1515
rect -1174 927 -1116 939
rect -716 1515 -658 1527
rect -716 939 -704 1515
rect -670 939 -658 1515
rect -716 927 -658 939
rect -258 1515 -200 1527
rect -258 939 -246 1515
rect -212 939 -200 1515
rect -258 927 -200 939
rect 200 1515 258 1527
rect 200 939 212 1515
rect 246 939 258 1515
rect 200 927 258 939
rect 658 1515 716 1527
rect 658 939 670 1515
rect 704 939 716 1515
rect 658 927 716 939
rect 1116 1515 1174 1527
rect 1116 939 1128 1515
rect 1162 939 1174 1515
rect 1116 927 1174 939
rect -1174 697 -1116 709
rect -1174 121 -1162 697
rect -1128 121 -1116 697
rect -1174 109 -1116 121
rect -716 697 -658 709
rect -716 121 -704 697
rect -670 121 -658 697
rect -716 109 -658 121
rect -258 697 -200 709
rect -258 121 -246 697
rect -212 121 -200 697
rect -258 109 -200 121
rect 200 697 258 709
rect 200 121 212 697
rect 246 121 258 697
rect 200 109 258 121
rect 658 697 716 709
rect 658 121 670 697
rect 704 121 716 697
rect 658 109 716 121
rect 1116 697 1174 709
rect 1116 121 1128 697
rect 1162 121 1174 697
rect 1116 109 1174 121
rect -1174 -121 -1116 -109
rect -1174 -697 -1162 -121
rect -1128 -697 -1116 -121
rect -1174 -709 -1116 -697
rect -716 -121 -658 -109
rect -716 -697 -704 -121
rect -670 -697 -658 -121
rect -716 -709 -658 -697
rect -258 -121 -200 -109
rect -258 -697 -246 -121
rect -212 -697 -200 -121
rect -258 -709 -200 -697
rect 200 -121 258 -109
rect 200 -697 212 -121
rect 246 -697 258 -121
rect 200 -709 258 -697
rect 658 -121 716 -109
rect 658 -697 670 -121
rect 704 -697 716 -121
rect 658 -709 716 -697
rect 1116 -121 1174 -109
rect 1116 -697 1128 -121
rect 1162 -697 1174 -121
rect 1116 -709 1174 -697
rect -1174 -939 -1116 -927
rect -1174 -1515 -1162 -939
rect -1128 -1515 -1116 -939
rect -1174 -1527 -1116 -1515
rect -716 -939 -658 -927
rect -716 -1515 -704 -939
rect -670 -1515 -658 -939
rect -716 -1527 -658 -1515
rect -258 -939 -200 -927
rect -258 -1515 -246 -939
rect -212 -1515 -200 -939
rect -258 -1527 -200 -1515
rect 200 -939 258 -927
rect 200 -1515 212 -939
rect 246 -1515 258 -939
rect 200 -1527 258 -1515
rect 658 -939 716 -927
rect 658 -1515 670 -939
rect 704 -1515 716 -939
rect 658 -1527 716 -1515
rect 1116 -939 1174 -927
rect 1116 -1515 1128 -939
rect 1162 -1515 1174 -939
rect 1116 -1527 1174 -1515
<< ndiffc >>
rect -1162 939 -1128 1515
rect -704 939 -670 1515
rect -246 939 -212 1515
rect 212 939 246 1515
rect 670 939 704 1515
rect 1128 939 1162 1515
rect -1162 121 -1128 697
rect -704 121 -670 697
rect -246 121 -212 697
rect 212 121 246 697
rect 670 121 704 697
rect 1128 121 1162 697
rect -1162 -697 -1128 -121
rect -704 -697 -670 -121
rect -246 -697 -212 -121
rect 212 -697 246 -121
rect 670 -697 704 -121
rect 1128 -697 1162 -121
rect -1162 -1515 -1128 -939
rect -704 -1515 -670 -939
rect -246 -1515 -212 -939
rect 212 -1515 246 -939
rect 670 -1515 704 -939
rect 1128 -1515 1162 -939
<< psubdiff >>
rect -1276 1667 -1180 1701
rect 1180 1667 1276 1701
rect -1276 1605 -1242 1667
rect 1242 1605 1276 1667
rect -1276 -1667 -1242 -1605
rect 1242 -1667 1276 -1605
rect -1276 -1701 -1180 -1667
rect 1180 -1701 1276 -1667
<< psubdiffcont >>
rect -1180 1667 1180 1701
rect -1276 -1605 -1242 1605
rect 1242 -1605 1276 1605
rect -1180 -1701 1180 -1667
<< poly >>
rect -1116 1599 -716 1615
rect -1116 1565 -1100 1599
rect -732 1565 -716 1599
rect -1116 1527 -716 1565
rect -658 1599 -258 1615
rect -658 1565 -642 1599
rect -274 1565 -258 1599
rect -658 1527 -258 1565
rect -200 1599 200 1615
rect -200 1565 -184 1599
rect 184 1565 200 1599
rect -200 1527 200 1565
rect 258 1599 658 1615
rect 258 1565 274 1599
rect 642 1565 658 1599
rect 258 1527 658 1565
rect 716 1599 1116 1615
rect 716 1565 732 1599
rect 1100 1565 1116 1599
rect 716 1527 1116 1565
rect -1116 889 -716 927
rect -1116 855 -1100 889
rect -732 855 -716 889
rect -1116 839 -716 855
rect -658 889 -258 927
rect -658 855 -642 889
rect -274 855 -258 889
rect -658 839 -258 855
rect -200 889 200 927
rect -200 855 -184 889
rect 184 855 200 889
rect -200 839 200 855
rect 258 889 658 927
rect 258 855 274 889
rect 642 855 658 889
rect 258 839 658 855
rect 716 889 1116 927
rect 716 855 732 889
rect 1100 855 1116 889
rect 716 839 1116 855
rect -1116 781 -716 797
rect -1116 747 -1100 781
rect -732 747 -716 781
rect -1116 709 -716 747
rect -658 781 -258 797
rect -658 747 -642 781
rect -274 747 -258 781
rect -658 709 -258 747
rect -200 781 200 797
rect -200 747 -184 781
rect 184 747 200 781
rect -200 709 200 747
rect 258 781 658 797
rect 258 747 274 781
rect 642 747 658 781
rect 258 709 658 747
rect 716 781 1116 797
rect 716 747 732 781
rect 1100 747 1116 781
rect 716 709 1116 747
rect -1116 71 -716 109
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 109
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 109
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 109
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -37 -716 -21
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -1116 -109 -716 -71
rect -658 -37 -258 -21
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -658 -109 -258 -71
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect 258 -37 658 -21
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 258 -109 658 -71
rect 716 -37 1116 -21
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 716 -109 1116 -71
rect -1116 -747 -716 -709
rect -1116 -781 -1100 -747
rect -732 -781 -716 -747
rect -1116 -797 -716 -781
rect -658 -747 -258 -709
rect -658 -781 -642 -747
rect -274 -781 -258 -747
rect -658 -797 -258 -781
rect -200 -747 200 -709
rect -200 -781 -184 -747
rect 184 -781 200 -747
rect -200 -797 200 -781
rect 258 -747 658 -709
rect 258 -781 274 -747
rect 642 -781 658 -747
rect 258 -797 658 -781
rect 716 -747 1116 -709
rect 716 -781 732 -747
rect 1100 -781 1116 -747
rect 716 -797 1116 -781
rect -1116 -855 -716 -839
rect -1116 -889 -1100 -855
rect -732 -889 -716 -855
rect -1116 -927 -716 -889
rect -658 -855 -258 -839
rect -658 -889 -642 -855
rect -274 -889 -258 -855
rect -658 -927 -258 -889
rect -200 -855 200 -839
rect -200 -889 -184 -855
rect 184 -889 200 -855
rect -200 -927 200 -889
rect 258 -855 658 -839
rect 258 -889 274 -855
rect 642 -889 658 -855
rect 258 -927 658 -889
rect 716 -855 1116 -839
rect 716 -889 732 -855
rect 1100 -889 1116 -855
rect 716 -927 1116 -889
rect -1116 -1565 -716 -1527
rect -1116 -1599 -1100 -1565
rect -732 -1599 -716 -1565
rect -1116 -1615 -716 -1599
rect -658 -1565 -258 -1527
rect -658 -1599 -642 -1565
rect -274 -1599 -258 -1565
rect -658 -1615 -258 -1599
rect -200 -1565 200 -1527
rect -200 -1599 -184 -1565
rect 184 -1599 200 -1565
rect -200 -1615 200 -1599
rect 258 -1565 658 -1527
rect 258 -1599 274 -1565
rect 642 -1599 658 -1565
rect 258 -1615 658 -1599
rect 716 -1565 1116 -1527
rect 716 -1599 732 -1565
rect 1100 -1599 1116 -1565
rect 716 -1615 1116 -1599
<< polycont >>
rect -1100 1565 -732 1599
rect -642 1565 -274 1599
rect -184 1565 184 1599
rect 274 1565 642 1599
rect 732 1565 1100 1599
rect -1100 855 -732 889
rect -642 855 -274 889
rect -184 855 184 889
rect 274 855 642 889
rect 732 855 1100 889
rect -1100 747 -732 781
rect -642 747 -274 781
rect -184 747 184 781
rect 274 747 642 781
rect 732 747 1100 781
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1100 -781 -732 -747
rect -642 -781 -274 -747
rect -184 -781 184 -747
rect 274 -781 642 -747
rect 732 -781 1100 -747
rect -1100 -889 -732 -855
rect -642 -889 -274 -855
rect -184 -889 184 -855
rect 274 -889 642 -855
rect 732 -889 1100 -855
rect -1100 -1599 -732 -1565
rect -642 -1599 -274 -1565
rect -184 -1599 184 -1565
rect 274 -1599 642 -1565
rect 732 -1599 1100 -1565
<< locali >>
rect -1276 1667 -1180 1701
rect 1180 1667 1276 1701
rect -1276 1605 -1242 1667
rect 1242 1605 1276 1667
rect -1116 1565 -1100 1599
rect -732 1565 -716 1599
rect -658 1565 -642 1599
rect -274 1565 -258 1599
rect -200 1565 -184 1599
rect 184 1565 200 1599
rect 258 1565 274 1599
rect 642 1565 658 1599
rect 716 1565 732 1599
rect 1100 1565 1116 1599
rect -1162 1515 -1128 1531
rect -1162 923 -1128 939
rect -704 1515 -670 1531
rect -704 923 -670 939
rect -246 1515 -212 1531
rect -246 923 -212 939
rect 212 1515 246 1531
rect 212 923 246 939
rect 670 1515 704 1531
rect 670 923 704 939
rect 1128 1515 1162 1531
rect 1128 923 1162 939
rect -1116 855 -1100 889
rect -732 855 -716 889
rect -658 855 -642 889
rect -274 855 -258 889
rect -200 855 -184 889
rect 184 855 200 889
rect 258 855 274 889
rect 642 855 658 889
rect 716 855 732 889
rect 1100 855 1116 889
rect -1116 747 -1100 781
rect -732 747 -716 781
rect -658 747 -642 781
rect -274 747 -258 781
rect -200 747 -184 781
rect 184 747 200 781
rect 258 747 274 781
rect 642 747 658 781
rect 716 747 732 781
rect 1100 747 1116 781
rect -1162 697 -1128 713
rect -1162 105 -1128 121
rect -704 697 -670 713
rect -704 105 -670 121
rect -246 697 -212 713
rect -246 105 -212 121
rect 212 697 246 713
rect 212 105 246 121
rect 670 697 704 713
rect 670 105 704 121
rect 1128 697 1162 713
rect 1128 105 1162 121
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect -1162 -121 -1128 -105
rect -1162 -713 -1128 -697
rect -704 -121 -670 -105
rect -704 -713 -670 -697
rect -246 -121 -212 -105
rect -246 -713 -212 -697
rect 212 -121 246 -105
rect 212 -713 246 -697
rect 670 -121 704 -105
rect 670 -713 704 -697
rect 1128 -121 1162 -105
rect 1128 -713 1162 -697
rect -1116 -781 -1100 -747
rect -732 -781 -716 -747
rect -658 -781 -642 -747
rect -274 -781 -258 -747
rect -200 -781 -184 -747
rect 184 -781 200 -747
rect 258 -781 274 -747
rect 642 -781 658 -747
rect 716 -781 732 -747
rect 1100 -781 1116 -747
rect -1116 -889 -1100 -855
rect -732 -889 -716 -855
rect -658 -889 -642 -855
rect -274 -889 -258 -855
rect -200 -889 -184 -855
rect 184 -889 200 -855
rect 258 -889 274 -855
rect 642 -889 658 -855
rect 716 -889 732 -855
rect 1100 -889 1116 -855
rect -1162 -939 -1128 -923
rect -1162 -1531 -1128 -1515
rect -704 -939 -670 -923
rect -704 -1531 -670 -1515
rect -246 -939 -212 -923
rect -246 -1531 -212 -1515
rect 212 -939 246 -923
rect 212 -1531 246 -1515
rect 670 -939 704 -923
rect 670 -1531 704 -1515
rect 1128 -939 1162 -923
rect 1128 -1531 1162 -1515
rect -1116 -1599 -1100 -1565
rect -732 -1599 -716 -1565
rect -658 -1599 -642 -1565
rect -274 -1599 -258 -1565
rect -200 -1599 -184 -1565
rect 184 -1599 200 -1565
rect 258 -1599 274 -1565
rect 642 -1599 658 -1565
rect 716 -1599 732 -1565
rect 1100 -1599 1116 -1565
rect -1276 -1667 -1242 -1605
rect 1242 -1667 1276 -1605
rect -1276 -1701 -1180 -1667
rect 1180 -1701 1276 -1667
<< viali >>
rect -1100 1565 -732 1599
rect -642 1565 -274 1599
rect -184 1565 184 1599
rect 274 1565 642 1599
rect 732 1565 1100 1599
rect -1162 939 -1128 1515
rect -704 939 -670 1515
rect -246 939 -212 1515
rect 212 939 246 1515
rect 670 939 704 1515
rect 1128 939 1162 1515
rect -1100 855 -732 889
rect -642 855 -274 889
rect -184 855 184 889
rect 274 855 642 889
rect 732 855 1100 889
rect -1100 747 -732 781
rect -642 747 -274 781
rect -184 747 184 781
rect 274 747 642 781
rect 732 747 1100 781
rect -1162 121 -1128 697
rect -704 121 -670 697
rect -246 121 -212 697
rect 212 121 246 697
rect 670 121 704 697
rect 1128 121 1162 697
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1162 -697 -1128 -121
rect -704 -697 -670 -121
rect -246 -697 -212 -121
rect 212 -697 246 -121
rect 670 -697 704 -121
rect 1128 -697 1162 -121
rect -1100 -781 -732 -747
rect -642 -781 -274 -747
rect -184 -781 184 -747
rect 274 -781 642 -747
rect 732 -781 1100 -747
rect -1100 -889 -732 -855
rect -642 -889 -274 -855
rect -184 -889 184 -855
rect 274 -889 642 -855
rect 732 -889 1100 -855
rect -1162 -1515 -1128 -939
rect -704 -1515 -670 -939
rect -246 -1515 -212 -939
rect 212 -1515 246 -939
rect 670 -1515 704 -939
rect 1128 -1515 1162 -939
rect -1100 -1599 -732 -1565
rect -642 -1599 -274 -1565
rect -184 -1599 184 -1565
rect 274 -1599 642 -1565
rect 732 -1599 1100 -1565
<< metal1 >>
rect -1112 1599 -720 1605
rect -1112 1565 -1100 1599
rect -732 1565 -720 1599
rect -1112 1559 -720 1565
rect -654 1599 -262 1605
rect -654 1565 -642 1599
rect -274 1565 -262 1599
rect -654 1559 -262 1565
rect -196 1599 196 1605
rect -196 1565 -184 1599
rect 184 1565 196 1599
rect -196 1559 196 1565
rect 262 1599 654 1605
rect 262 1565 274 1599
rect 642 1565 654 1599
rect 262 1559 654 1565
rect 720 1599 1112 1605
rect 720 1565 732 1599
rect 1100 1565 1112 1599
rect 720 1559 1112 1565
rect -1168 1515 -1122 1527
rect -1168 939 -1162 1515
rect -1128 939 -1122 1515
rect -1168 927 -1122 939
rect -710 1515 -664 1527
rect -710 939 -704 1515
rect -670 939 -664 1515
rect -710 927 -664 939
rect -252 1515 -206 1527
rect -252 939 -246 1515
rect -212 939 -206 1515
rect -252 927 -206 939
rect 206 1515 252 1527
rect 206 939 212 1515
rect 246 939 252 1515
rect 206 927 252 939
rect 664 1515 710 1527
rect 664 939 670 1515
rect 704 939 710 1515
rect 664 927 710 939
rect 1122 1515 1168 1527
rect 1122 939 1128 1515
rect 1162 939 1168 1515
rect 1122 927 1168 939
rect -1112 889 -720 895
rect -1112 855 -1100 889
rect -732 855 -720 889
rect -1112 849 -720 855
rect -654 889 -262 895
rect -654 855 -642 889
rect -274 855 -262 889
rect -654 849 -262 855
rect -196 889 196 895
rect -196 855 -184 889
rect 184 855 196 889
rect -196 849 196 855
rect 262 889 654 895
rect 262 855 274 889
rect 642 855 654 889
rect 262 849 654 855
rect 720 889 1112 895
rect 720 855 732 889
rect 1100 855 1112 889
rect 720 849 1112 855
rect -1112 781 -720 787
rect -1112 747 -1100 781
rect -732 747 -720 781
rect -1112 741 -720 747
rect -654 781 -262 787
rect -654 747 -642 781
rect -274 747 -262 781
rect -654 741 -262 747
rect -196 781 196 787
rect -196 747 -184 781
rect 184 747 196 781
rect -196 741 196 747
rect 262 781 654 787
rect 262 747 274 781
rect 642 747 654 781
rect 262 741 654 747
rect 720 781 1112 787
rect 720 747 732 781
rect 1100 747 1112 781
rect 720 741 1112 747
rect -1168 697 -1122 709
rect -1168 121 -1162 697
rect -1128 121 -1122 697
rect -1168 109 -1122 121
rect -710 697 -664 709
rect -710 121 -704 697
rect -670 121 -664 697
rect -710 109 -664 121
rect -252 697 -206 709
rect -252 121 -246 697
rect -212 121 -206 697
rect -252 109 -206 121
rect 206 697 252 709
rect 206 121 212 697
rect 246 121 252 697
rect 206 109 252 121
rect 664 697 710 709
rect 664 121 670 697
rect 704 121 710 697
rect 664 109 710 121
rect 1122 697 1168 709
rect 1122 121 1128 697
rect 1162 121 1168 697
rect 1122 109 1168 121
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1112 -37 -720 -31
rect -1112 -71 -1100 -37
rect -732 -71 -720 -37
rect -1112 -77 -720 -71
rect -654 -37 -262 -31
rect -654 -71 -642 -37
rect -274 -71 -262 -37
rect -654 -77 -262 -71
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect 262 -37 654 -31
rect 262 -71 274 -37
rect 642 -71 654 -37
rect 262 -77 654 -71
rect 720 -37 1112 -31
rect 720 -71 732 -37
rect 1100 -71 1112 -37
rect 720 -77 1112 -71
rect -1168 -121 -1122 -109
rect -1168 -697 -1162 -121
rect -1128 -697 -1122 -121
rect -1168 -709 -1122 -697
rect -710 -121 -664 -109
rect -710 -697 -704 -121
rect -670 -697 -664 -121
rect -710 -709 -664 -697
rect -252 -121 -206 -109
rect -252 -697 -246 -121
rect -212 -697 -206 -121
rect -252 -709 -206 -697
rect 206 -121 252 -109
rect 206 -697 212 -121
rect 246 -697 252 -121
rect 206 -709 252 -697
rect 664 -121 710 -109
rect 664 -697 670 -121
rect 704 -697 710 -121
rect 664 -709 710 -697
rect 1122 -121 1168 -109
rect 1122 -697 1128 -121
rect 1162 -697 1168 -121
rect 1122 -709 1168 -697
rect -1112 -747 -720 -741
rect -1112 -781 -1100 -747
rect -732 -781 -720 -747
rect -1112 -787 -720 -781
rect -654 -747 -262 -741
rect -654 -781 -642 -747
rect -274 -781 -262 -747
rect -654 -787 -262 -781
rect -196 -747 196 -741
rect -196 -781 -184 -747
rect 184 -781 196 -747
rect -196 -787 196 -781
rect 262 -747 654 -741
rect 262 -781 274 -747
rect 642 -781 654 -747
rect 262 -787 654 -781
rect 720 -747 1112 -741
rect 720 -781 732 -747
rect 1100 -781 1112 -747
rect 720 -787 1112 -781
rect -1112 -855 -720 -849
rect -1112 -889 -1100 -855
rect -732 -889 -720 -855
rect -1112 -895 -720 -889
rect -654 -855 -262 -849
rect -654 -889 -642 -855
rect -274 -889 -262 -855
rect -654 -895 -262 -889
rect -196 -855 196 -849
rect -196 -889 -184 -855
rect 184 -889 196 -855
rect -196 -895 196 -889
rect 262 -855 654 -849
rect 262 -889 274 -855
rect 642 -889 654 -855
rect 262 -895 654 -889
rect 720 -855 1112 -849
rect 720 -889 732 -855
rect 1100 -889 1112 -855
rect 720 -895 1112 -889
rect -1168 -939 -1122 -927
rect -1168 -1515 -1162 -939
rect -1128 -1515 -1122 -939
rect -1168 -1527 -1122 -1515
rect -710 -939 -664 -927
rect -710 -1515 -704 -939
rect -670 -1515 -664 -939
rect -710 -1527 -664 -1515
rect -252 -939 -206 -927
rect -252 -1515 -246 -939
rect -212 -1515 -206 -939
rect -252 -1527 -206 -1515
rect 206 -939 252 -927
rect 206 -1515 212 -939
rect 246 -1515 252 -939
rect 206 -1527 252 -1515
rect 664 -939 710 -927
rect 664 -1515 670 -939
rect 704 -1515 710 -939
rect 664 -1527 710 -1515
rect 1122 -939 1168 -927
rect 1122 -1515 1128 -939
rect 1162 -1515 1168 -939
rect 1122 -1527 1168 -1515
rect -1112 -1565 -720 -1559
rect -1112 -1599 -1100 -1565
rect -732 -1599 -720 -1565
rect -1112 -1605 -720 -1599
rect -654 -1565 -262 -1559
rect -654 -1599 -642 -1565
rect -274 -1599 -262 -1565
rect -654 -1605 -262 -1599
rect -196 -1565 196 -1559
rect -196 -1599 -184 -1565
rect 184 -1599 196 -1565
rect -196 -1605 196 -1599
rect 262 -1565 654 -1559
rect 262 -1599 274 -1565
rect 642 -1599 654 -1565
rect 262 -1605 654 -1599
rect 720 -1565 1112 -1559
rect 720 -1599 732 -1565
rect 1100 -1599 1112 -1565
rect 720 -1605 1112 -1599
<< properties >>
string FIXED_BBOX -1259 -1684 1259 1684
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 2.0 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
