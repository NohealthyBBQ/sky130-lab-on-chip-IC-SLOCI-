magic
tech sky130A
magscale 1 2
timestamp 1662486269
<< pwell >>
rect -307 -2198 307 2198
<< psubdiff >>
rect -271 2128 -175 2162
rect 175 2128 271 2162
rect -271 2066 -237 2128
rect 237 2066 271 2128
rect -271 -2128 -237 -2066
rect 237 -2128 271 -2066
rect -271 -2162 -175 -2128
rect 175 -2162 271 -2128
<< psubdiffcont >>
rect -175 2128 175 2162
rect -271 -2066 -237 2066
rect 237 -2066 271 2066
rect -175 -2162 175 -2128
<< xpolycontact >>
rect -141 1600 141 2032
rect -141 -2032 141 -1600
<< ppolyres >>
rect -141 -1600 141 1600
<< locali >>
rect -271 2128 -175 2162
rect 175 2128 271 2162
rect -271 2066 -237 2128
rect 237 2066 271 2128
rect -271 -2128 -237 -2066
rect 237 -2128 271 -2066
rect -271 -2162 -175 -2128
rect 175 -2162 271 -2128
<< viali >>
rect -125 1617 125 2014
rect -125 -2014 125 -1617
<< metal1 >>
rect -131 2014 131 2026
rect -131 1617 -125 2014
rect 125 1617 131 2014
rect -131 1605 131 1617
rect -131 -1617 131 -1605
rect -131 -2014 -125 -1617
rect 125 -2014 131 -1617
rect -131 -2026 131 -2014
<< res1p41 >>
rect -143 -1602 143 1602
<< properties >>
string FIXED_BBOX -254 -2145 254 2145
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 16.0 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 3.905k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
