magic
tech sky130A
magscale 1 2
timestamp 1661869741
<< metal1 >>
rect 522 2926 532 3026
rect 612 2926 622 3026
rect 1438 2926 1448 3026
rect 1528 2926 1538 3026
rect 2352 2926 2362 3026
rect 2442 2926 2452 3026
rect 1465 2916 1471 2926
rect 1505 2916 1511 2926
rect 2379 2916 2385 2926
rect 2419 2916 2425 2926
rect 1921 2536 1927 2546
rect 1961 2536 1967 2546
rect 1007 2524 1013 2534
rect 1047 2524 1053 2534
rect 64 2424 74 2524
rect 154 2424 164 2524
rect 980 2424 990 2524
rect 1070 2424 1080 2524
rect 1894 2436 1904 2536
rect 1984 2436 1994 2536
rect 527 2347 617 2393
rect 985 2347 1075 2393
rect 1443 2347 1533 2393
rect 1901 2347 1991 2393
rect 89 2257 135 2269
rect 89 1768 95 2257
rect 129 1768 135 2257
rect 520 2170 530 2270
rect 610 2170 620 2270
rect 1005 2257 1051 2269
rect 62 1668 72 1768
rect 152 1668 162 1768
rect 547 1681 553 2170
rect 587 1681 593 2170
rect 1005 1768 1011 2257
rect 1045 1768 1051 2257
rect 1436 2170 1446 2270
rect 1526 2170 1536 2270
rect 1921 2257 1967 2269
rect 547 1669 593 1681
rect 978 1668 988 1768
rect 1068 1668 1078 1768
rect 1463 1681 1469 2170
rect 1503 1681 1509 2170
rect 1921 1790 1927 2257
rect 1961 1790 1967 2257
rect 2350 2170 2360 2270
rect 2440 2170 2450 2270
rect 2377 2160 2385 2170
rect 2417 2160 2425 2170
rect 1919 1780 1927 1790
rect 1959 1780 1967 1790
rect 1463 1669 1509 1681
rect 1892 1680 1902 1780
rect 1982 1680 1992 1780
rect 2379 1681 2385 2160
rect 2419 1681 2425 2160
rect 1921 1669 1967 1680
rect 2379 1669 2425 1681
rect 527 1591 617 1637
rect 985 1591 1075 1637
rect 1443 1591 1533 1637
rect 1901 1591 1991 1637
rect 91 1501 137 1513
rect 91 1012 97 1501
rect 131 1012 137 1501
rect 522 1414 532 1514
rect 612 1414 622 1514
rect 1007 1501 1053 1513
rect 64 912 74 1012
rect 154 912 164 1012
rect 549 925 555 1414
rect 589 925 595 1414
rect 1007 1012 1013 1501
rect 1047 1012 1053 1501
rect 1438 1414 1448 1514
rect 1528 1414 1538 1514
rect 1923 1501 1969 1513
rect 549 913 595 925
rect 980 912 990 1012
rect 1070 912 1080 1012
rect 1465 925 1471 1414
rect 1505 925 1511 1414
rect 1923 1034 1929 1501
rect 1963 1034 1969 1501
rect 2352 1414 2362 1514
rect 2442 1414 2452 1514
rect 2379 1404 2387 1414
rect 2419 1404 2427 1414
rect 1921 1024 1929 1034
rect 1961 1024 1969 1034
rect 1465 913 1511 925
rect 1894 924 1904 1024
rect 1984 924 1994 1024
rect 2381 925 2387 1404
rect 2421 925 2427 1404
rect 1923 913 1969 924
rect 2381 913 2427 925
rect 527 835 617 881
rect 985 835 1075 881
rect 1443 835 1533 881
rect 1901 835 1991 881
rect 91 745 137 757
rect 91 256 97 745
rect 131 256 137 745
rect 522 658 532 758
rect 612 658 622 758
rect 1007 745 1053 757
rect 64 156 74 256
rect 154 156 164 256
rect 549 169 555 658
rect 589 169 595 658
rect 1007 256 1013 745
rect 1047 256 1053 745
rect 1438 658 1448 758
rect 1528 658 1538 758
rect 1923 745 1969 757
rect 549 157 595 169
rect 980 156 990 256
rect 1070 156 1080 256
rect 1465 169 1471 658
rect 1505 169 1511 658
rect 1923 278 1929 745
rect 1963 278 1969 745
rect 2352 658 2362 758
rect 2442 658 2452 758
rect 2379 648 2387 658
rect 2419 648 2427 658
rect 1921 268 1929 278
rect 1961 268 1969 278
rect 1465 157 1511 169
rect 1894 168 1904 268
rect 1984 168 1994 268
rect 2381 169 2387 648
rect 2421 169 2427 648
rect 1923 157 1969 168
rect 2381 157 2427 169
rect 527 79 617 125
rect 985 79 1075 125
rect 1443 79 1533 125
rect 1901 79 1991 125
<< via1 >>
rect 532 2926 612 3026
rect 1448 2926 1528 3026
rect 2362 2926 2442 3026
rect 74 2424 154 2524
rect 990 2424 1070 2524
rect 1904 2436 1984 2536
rect 530 2170 610 2270
rect 72 1668 152 1768
rect 1446 2170 1526 2270
rect 988 1668 1068 1768
rect 2360 2170 2440 2270
rect 1902 1680 1982 1780
rect 532 1414 612 1514
rect 74 912 154 1012
rect 1448 1414 1528 1514
rect 990 912 1070 1012
rect 2362 1414 2442 1514
rect 1904 924 1984 1024
rect 532 658 612 758
rect 74 156 154 256
rect 1448 658 1528 758
rect 990 156 1070 256
rect 2362 658 2442 758
rect 1904 168 1984 268
<< metal2 >>
rect 532 3026 612 3036
rect 532 2916 612 2926
rect 1448 3026 1528 3036
rect 1448 2916 1528 2926
rect 2362 3026 2442 3036
rect 2362 2916 2442 2926
rect 1904 2536 1984 2546
rect 74 2524 154 2534
rect 74 2414 154 2424
rect 990 2524 1070 2534
rect 1904 2426 1984 2436
rect 990 2414 1070 2424
rect 530 2270 610 2280
rect 530 2160 610 2170
rect 1446 2270 1526 2280
rect 1446 2160 1526 2170
rect 2360 2270 2440 2280
rect 2360 2160 2440 2170
rect 1902 1780 1982 1790
rect 72 1768 152 1778
rect 72 1658 152 1668
rect 988 1768 1068 1778
rect 1902 1670 1982 1680
rect 988 1658 1068 1668
rect 532 1514 612 1524
rect 532 1404 612 1414
rect 1448 1514 1528 1524
rect 1448 1404 1528 1414
rect 2362 1514 2442 1524
rect 2362 1404 2442 1414
rect 1904 1024 1984 1034
rect 74 1012 154 1022
rect 74 902 154 912
rect 990 1012 1070 1022
rect 1904 914 1984 924
rect 990 902 1070 912
rect 532 758 612 768
rect 532 648 612 658
rect 1448 758 1528 768
rect 1448 648 1528 658
rect 2362 758 2442 768
rect 2362 648 2442 658
rect 1904 268 1984 278
rect 74 256 154 266
rect 74 146 154 156
rect 990 256 1070 266
rect 1904 158 1984 168
rect 990 146 1070 156
use sky130_fd_pr__nfet_01v8_USQY94  sky130_fd_pr__nfet_01v8_USQY94_0
timestamp 1661796674
transform 1 0 1259 0 1 1560
box -1312 -1613 1312 1613
<< end >>
