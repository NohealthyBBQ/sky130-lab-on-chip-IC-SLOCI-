magic
tech sky130A
magscale 1 2
timestamp 1661816812
<< metal1 >>
rect 527 2347 617 2393
rect 985 2353 1075 2387
rect 1443 2347 1533 2393
rect 1901 2347 1991 2393
rect 527 1591 617 1637
rect 985 1591 1075 1637
rect 1443 1591 1533 1637
rect 1901 1591 1991 1637
rect 527 835 617 881
rect 985 835 1075 881
rect 1443 835 1533 881
rect 1901 835 1991 881
rect 985 79 1075 125
rect 1443 79 1533 125
rect 1901 79 1991 125
use sky130_fd_pr__nfet_01v8_USQY94  sky130_fd_pr__nfet_01v8_USQY94_0
timestamp 1661796674
transform 1 0 1259 0 1 1560
box -1312 -1613 1312 1613
<< end >>
